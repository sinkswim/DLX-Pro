
module DLX ( clk, rst, iram_data, Data_out_fromRAM, addr_to_iram, read_op, 
        write_op, nibble, write_byte, Address_toRAM, Data_in );
  input [31:0] iram_data;
  input [31:0] Data_out_fromRAM;
  output [31:0] addr_to_iram;
  output [1:0] nibble;
  output [31:0] Address_toRAM;
  output [31:0] Data_in;
  input clk, rst;
  output read_op, write_op, write_byte;
  wire   n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, \u_DataPath/reg_write_i ,
         \u_DataPath/jump_i , \u_DataPath/u_fetch/pc1/N3 ,
         \u_DataPath/u_decode_unit/reg_file0/N154 ,
         \u_DataPath/u_decode_unit/reg_file0/N153 ,
         \u_DataPath/u_decode_unit/reg_file0/N152 ,
         \u_DataPath/u_decode_unit/reg_file0/N151 ,
         \u_DataPath/u_decode_unit/reg_file0/N150 ,
         \u_DataPath/u_decode_unit/reg_file0/N149 ,
         \u_DataPath/u_decode_unit/reg_file0/N148 ,
         \u_DataPath/u_decode_unit/reg_file0/N147 ,
         \u_DataPath/u_decode_unit/reg_file0/N146 ,
         \u_DataPath/u_decode_unit/reg_file0/N145 ,
         \u_DataPath/u_decode_unit/reg_file0/N144 ,
         \u_DataPath/u_decode_unit/reg_file0/N143 ,
         \u_DataPath/u_decode_unit/reg_file0/N142 ,
         \u_DataPath/u_decode_unit/reg_file0/N141 ,
         \u_DataPath/u_decode_unit/reg_file0/N140 ,
         \u_DataPath/u_decode_unit/reg_file0/N139 ,
         \u_DataPath/u_decode_unit/reg_file0/N138 ,
         \u_DataPath/u_decode_unit/reg_file0/N137 ,
         \u_DataPath/u_decode_unit/reg_file0/N136 ,
         \u_DataPath/u_decode_unit/reg_file0/N135 ,
         \u_DataPath/u_decode_unit/reg_file0/N134 ,
         \u_DataPath/u_decode_unit/reg_file0/N133 ,
         \u_DataPath/u_decode_unit/reg_file0/N132 ,
         \u_DataPath/u_decode_unit/reg_file0/N131 ,
         \u_DataPath/u_decode_unit/reg_file0/N130 ,
         \u_DataPath/u_decode_unit/reg_file0/N129 ,
         \u_DataPath/u_decode_unit/reg_file0/N128 ,
         \u_DataPath/u_decode_unit/reg_file0/N127 ,
         \u_DataPath/u_decode_unit/reg_file0/N126 ,
         \u_DataPath/u_decode_unit/reg_file0/N125 ,
         \u_DataPath/u_decode_unit/reg_file0/N92 ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ,
         \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ,
         \u_DataPath/u_idexreg/N184 , \u_DataPath/u_idexreg/N33 ,
         \u_DataPath/u_idexreg/N31 , \u_DataPath/u_idexreg/N16 ,
         \u_DataPath/u_idexreg/N15 , \u_DataPath/u_idexreg/N10 ,
         \u_DataPath/u_idexreg/N3 , \u_DataPath/u_execute/ovf_i ,
         \u_DataPath/u_execute/EXALU/N811 , \u_DataPath/u_execute/EXALU/N810 ,
         \u_DataPath/u_exmemreg/N78 , \u_DataPath/u_memwbreg/N64 , n2733,
         \lte_x_59/B[28] , \lte_x_59/B[26] , \lte_x_59/B[24] ,
         \lte_x_59/B[22] , \lte_x_59/B[21] , \lte_x_59/B[18] ,
         \lte_x_59/B[16] , \lte_x_59/B[15] , \lte_x_59/B[14] , \lte_x_59/B[9] ,
         \lte_x_59/B[8] , \lte_x_59/B[7] , \lte_x_59/B[6] , \lte_x_59/B[5] ,
         \lte_x_59/B[4] , \lte_x_59/B[3] , \lte_x_59/B[1] , \sub_x_53/A[30] ,
         \sub_x_53/A[29] , \sub_x_53/A[27] , \sub_x_53/A[25] ,
         \sub_x_53/A[23] , \sub_x_53/A[20] , \sub_x_53/A[17] , \sub_x_53/A[2] ,
         \sub_x_53/A[0] , n2773, n2774, n2776, n2778, n2780, n2782, n2784,
         n2787, n2789, n2791, n2793, n2795, n2797, n2799, n2801, n2803, n2805,
         n2807, n2809, n2811, n2813, n2815, n2817, n2819, n2821, n2823, n2825,
         n2829, n2831, n2833, n2835, n2838, n2840, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2851, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2864, n2865, n2866, n2867, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2993, n2994, n2995, n2996,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3018,
         n3020, n3021, n3022, n3023, n3024, n3025, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3066, n3067, n3068, n3069, n3070, n3072, n3073, n3074,
         n3075, n3076, n3077, n3079, n3080, n3081, n3082, n3084, n3085, n3086,
         n3088, n3089, n3090, n3091, n3093, n3094, n3095, n3096, n3098, n3099,
         n3100, n3101, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4823, n4824, n4825, n4826, n4827, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5224, n5225, n5226, n5227, n5228, n5229, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5777, n5778, n5779, n5780, n5781, n5782, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5841, n5842, n5844, n5845, n5846, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5989, n5990, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6034, n6035, n6036, n6037, n6038, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6087, n6088, n6089, n6090, n6091, n6092,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7652, n7653, n7654, n7655, n7657, n7658, n7659,
         n7660, n7661, n7663, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7676, n7677, n7678, n7679, n7680, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7749, n7750, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7877, n7878, n7879, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7913, n7914, n7915, n7916, n7917, n7918, n7920, n7921, n7922,
         n7923, n7924, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8190, n8191, n8193, n8194, n8196, n8197, n8198,
         n8200, n8202, n8204, n8205, n8206, n8208, n8209, n8211, n8212, n8213,
         n8214, n8216, n8218, n8219, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8233, n8234, n8235, n8236, n8238,
         n8240, n8242, n8243, n8245, n8247, n8251, n8253, n8255, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8277, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8585, n8586,
         n8587, n8588, n8589, n8591, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8616, n8618, n8620, n8621,
         n8622, n8623, n8625, n8626, n8627, n8629, n8631, n8634, n8635, n8636,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9352, n9354, n9355, n9356, n9357, n9359, n9360,
         n9361, n9362, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9431;
  wire   [5:0] opcode_i;
  wire   [4:0] \u_DataPath/regfile_addr_out_towb_i ;
  wire   [31:0] \u_DataPath/from_alu_data_out_i ;
  wire   [31:0] \u_DataPath/from_mem_data_out_i ;
  wire   [2:0] \u_DataPath/cw_towb_i ;
  wire   [4:0] \u_DataPath/RFaddr_out_memwb_i ;
  wire   [31:0] \u_DataPath/dataOut_exe_i ;
  wire   [2:0] \u_DataPath/cw_memwb_i ;
  wire   [31:0] \u_DataPath/mem_writedata_out_i ;
  wire   [10:0] \u_DataPath/cw_tomem_i ;
  wire   [31:0] \u_DataPath/toPC2_i ;
  wire   [10:0] \u_DataPath/cw_exmem_i ;
  wire   [4:0] \u_DataPath/rs_ex_i ;
  wire   [31:0] \u_DataPath/immediate_ext_ex_i ;
  wire   [31:0] \u_DataPath/data_read_ex_2_i ;
  wire   [31:0] \u_DataPath/data_read_ex_1_i ;
  wire   [31:0] \u_DataPath/pc_4_to_ex_i ;
  wire   [21:0] \u_DataPath/cw_to_ex_i ;
  wire   [31:0] \u_DataPath/immediate_ext_dec_i ;
  wire   [31:0] \u_DataPath/pc4_to_idexreg_i ;
  wire   [31:0] \u_DataPath/jaddr_i ;
  wire   [4:0] \u_DataPath/idex_rt_i ;
  wire   [31:0] \u_DataPath/pc_4_i ;
  wire   [31:0] \u_DataPath/branch_target_i ;
  wire   [31:0] \u_DataPath/jump_address_i ;
  wire   [1:0] \u_DataPath/u_decode_unit/hdu_0/current_state ;
  wire   [31:0] \u_DataPath/u_execute/psw_status_i ;
  wire   [31:0] \u_DataPath/u_execute/link_value_i ;
  wire   [31:0] \u_DataPath/u_execute/resAdd1_i ;
  assign Address_toRAM[30] = 1'b0;
  assign Address_toRAM[31] = 1'b0;
  assign addr_to_iram[30] = 1'b0;
  assign addr_to_iram[31] = 1'b0;

  HS65_LH_CNIVX3 U151 ( .A(rst), .Z(n2733) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[19][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N136 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[4][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N151 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[5][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N150 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_execute/EXALU/ovf_reg  ( .G(
        \u_DataPath/u_execute/EXALU/N810 ), .D(
        \u_DataPath/u_execute/EXALU/N811 ), .Q(\u_DataPath/u_execute/ovf_i )
         );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[3][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N152 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[9][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N146 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[17][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N138 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[27][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N128 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[25][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N130 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[13][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N142 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[11][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N144 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[10][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N145 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[1][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N154 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[20][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N135 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[2][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N153 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[6][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N149 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[15][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N140 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[12][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N143 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[16][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N139 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[8][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N147 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[24][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N131 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8030), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n8021), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[14][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N141 ), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[21][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N134 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7999), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8026), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8017), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][6]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8016), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7981), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7936), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][2]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8029), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7954), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][16]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7953), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7960), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7938), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8032), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7978), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8014), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7993), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][25]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7992), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8023), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][5]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8022), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8008), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][29]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8007), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7951), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7969), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7996), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8005), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7945), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][10]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7944), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7962), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7942), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7972), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][15]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7971), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[22][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N133 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][31]  ( 
        .G(rst), .D(n7937), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][0]  ( 
        .G(rst), .D(n8000), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][1]  ( 
        .G(rst), .D(n8027), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][6]  ( 
        .G(rst), .D(n8018), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][18]  ( 
        .G(rst), .D(n7982), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][2]  ( 
        .G(rst), .D(n8028), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][17]  ( 
        .G(rst), .D(n7988), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][16]  ( 
        .G(rst), .D(n7955), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][20]  ( 
        .G(rst), .D(n7961), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][8]  ( 
        .G(rst), .D(n7940), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][4]  ( 
        .G(rst), .D(n8033), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][22]  ( 
        .G(rst), .D(n7979), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][28]  ( 
        .G(rst), .D(n7931), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][24]  ( 
        .G(rst), .D(n7985), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][9]  ( 
        .G(rst), .D(n8015), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][25]  ( 
        .G(rst), .D(n7994), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][5]  ( 
        .G(rst), .D(n8024), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][21]  ( 
        .G(rst), .D(n7967), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][29]  ( 
        .G(rst), .D(n8009), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][13]  ( 
        .G(rst), .D(n7958), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][7]  ( 
        .G(rst), .D(n7952), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][12]  ( 
        .G(rst), .D(n7970), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][30]  ( 
        .G(rst), .D(n8011), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][23]  ( 
        .G(rst), .D(n7997), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][26]  ( 
        .G(rst), .D(n8006), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][10]  ( 
        .G(rst), .D(n7946), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][3]  ( 
        .G(rst), .D(n8020), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][19]  ( 
        .G(rst), .D(n7964), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][11]  ( 
        .G(rst), .D(n7943), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][15]  ( 
        .G(rst), .D(n7973), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][14]  ( 
        .G(rst), .D(n7991), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[0][27]  ( 
        .G(rst), .D(n7928), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ) );
  HS65_LH_LDHQX9 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[7][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N148 ), .D(n8010), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][31]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7935), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][26]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n8004), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7930), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][19]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7963), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[23][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N132 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][18]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7980), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][4]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8031), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][3]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8019), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][1]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8025), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7966), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7927), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ) );
  HS65_LL_IVX18 U3438 ( .A(n3118), .Z(addr_to_iram[26]) );
  HS65_LH_IVX40 U3462 ( .A(n2782), .Z(addr_to_iram[17]) );
  HS65_LH_IVX40 U3463 ( .A(n2823), .Z(addr_to_iram[9]) );
  HS65_LH_IVX40 U3464 ( .A(n2825), .Z(addr_to_iram[25]) );
  HS65_LH_IVX40 U3466 ( .A(n2829), .Z(addr_to_iram[7]) );
  HS65_LH_IVX40 U3467 ( .A(n2831), .Z(addr_to_iram[18]) );
  HS65_LH_IVX40 U3468 ( .A(n2833), .Z(addr_to_iram[8]) );
  HS65_LH_IVX40 U3469 ( .A(n2835), .Z(addr_to_iram[6]) );
  HS65_LH_NOR4ABX2 U3470 ( .A(n6806), .B(n6805), .C(n6804), .D(n6803), .Z(
        n8183) );
  HS65_LH_NOR4ABX2 U3471 ( .A(n6846), .B(n6845), .C(n6844), .D(n6843), .Z(
        n8156) );
  HS65_LL_OR2ABX35 U3473 ( .A(n2981), .B(n2994), .Z(write_op) );
  HS65_LH_IVX9 U3474 ( .A(n3003), .Z(n2787) );
  HS65_LH_IVX9 U3475 ( .A(n3004), .Z(n2793) );
  HS65_LH_IVX9 U3476 ( .A(n2993), .Z(n2809) );
  HS65_LH_IVX9 U3477 ( .A(n3006), .Z(n2805) );
  HS65_LH_IVX9 U3478 ( .A(n3005), .Z(n2803) );
  HS65_LH_IVX9 U3479 ( .A(n3007), .Z(n2807) );
  HS65_LH_IVX9 U3480 ( .A(n8687), .Z(\u_DataPath/pc_4_i [2]) );
  HS65_LH_IVX9 U3481 ( .A(n2989), .Z(n2789) );
  HS65_LH_IVX9 U3482 ( .A(n2987), .Z(n2791) );
  HS65_LH_IVX9 U3483 ( .A(n3001), .Z(n2795) );
  HS65_LH_IVX9 U3484 ( .A(n3000), .Z(n2797) );
  HS65_LH_IVX9 U3485 ( .A(n3002), .Z(n2799) );
  HS65_LH_IVX9 U3486 ( .A(n2996), .Z(n2813) );
  HS65_LH_IVX9 U3487 ( .A(n2999), .Z(n2815) );
  HS65_LH_IVX9 U3488 ( .A(n2995), .Z(n2817) );
  HS65_LH_IVX9 U3489 ( .A(n8671), .Z(n2774) );
  HS65_LH_IVX9 U3490 ( .A(n8675), .Z(n2776) );
  HS65_LH_IVX9 U3491 ( .A(n8673), .Z(n2778) );
  HS65_LH_IVX9 U3492 ( .A(n8672), .Z(n2819) );
  HS65_LH_IVX9 U3493 ( .A(n8674), .Z(n2821) );
  HS65_LH_IVX9 U3494 ( .A(n3013), .Z(n2838) );
  HS65_LH_IVX9 U3495 ( .A(n2998), .Z(n2811) );
  HS65_LH_IVX9 U3496 ( .A(n8692), .Z(n2782) );
  HS65_LH_IVX9 U3497 ( .A(n8703), .Z(n2825) );
  HS65_LH_IVX9 U3498 ( .A(n8679), .Z(n2823) );
  HS65_LH_IVX9 U3500 ( .A(n8678), .Z(n2829) );
  HS65_LH_IVX9 U3501 ( .A(n8697), .Z(n2831) );
  HS65_LH_IVX9 U3502 ( .A(n8681), .Z(n2833) );
  HS65_LH_IVX9 U3503 ( .A(n8680), .Z(n2835) );
  HS65_LH_IVX9 U3504 ( .A(n8684), .Z(n7745) );
  HS65_LH_IVX9 U3505 ( .A(n8686), .Z(n3126) );
  HS65_LH_IVX9 U3506 ( .A(n8685), .Z(n7669) );
  HS65_LH_AOI21X2 U3507 ( .A(n7631), .B(n5707), .C(n5706), .Z(n5709) );
  HS65_LH_NOR2AX3 U3517 ( .A(\u_DataPath/dataOut_exe_i [29]), .B(n3116), .Z(
        n2988) );
  HS65_LH_NOR2AX3 U3518 ( .A(n8748), .B(n3115), .Z(n2998) );
  HS65_LH_AOI21X2 U3519 ( .A(n6011), .B(n6083), .C(n6010), .Z(n6065) );
  HS65_LH_IVX9 U3520 ( .A(n8713), .Z(n2780) );
  HS65_LH_AOI21X2 U3521 ( .A(n6117), .B(n6119), .C(n5943), .Z(n2876) );
  HS65_LL_NAND3AX6 U3522 ( .A(n5676), .B(n8478), .C(n5675), .Z(n5677) );
  HS65_LH_BFX9 U3523 ( .A(n7096), .Z(n7902) );
  HS65_LH_BFX9 U3528 ( .A(n7320), .Z(n7587) );
  HS65_LH_BFX9 U3529 ( .A(n7330), .Z(n7600) );
  HS65_LH_BFX9 U3530 ( .A(n7332), .Z(n7602) );
  HS65_LH_BFX9 U3531 ( .A(n7317), .Z(n7585) );
  HS65_LH_BFX9 U3532 ( .A(n6675), .Z(n7318) );
  HS65_LH_BFX9 U3533 ( .A(n7311), .Z(n7579) );
  HS65_LH_AOI21X2 U3534 ( .A(Data_out_fromRAM[15]), .B(n8271), .C(n7344), .Z(
        n7345) );
  HS65_LH_BFX9 U3535 ( .A(n6382), .Z(n7291) );
  HS65_LH_BFX9 U3537 ( .A(n6681), .Z(n7523) );
  HS65_LH_NOR2X6 U3541 ( .A(n6348), .B(n2878), .Z(n7578) );
  HS65_LH_NOR2X6 U3542 ( .A(n6147), .B(n6153), .Z(n6617) );
  HS65_LH_NOR2X6 U3543 ( .A(n6150), .B(n6147), .Z(n6162) );
  HS65_LH_NOR2X6 U3545 ( .A(n6153), .B(n6140), .Z(n6635) );
  HS65_LH_NOR2X6 U3546 ( .A(n6353), .B(n6352), .Z(n6967) );
  HS65_LH_NOR2X6 U3548 ( .A(n6349), .B(n6332), .Z(n7311) );
  HS65_LH_NOR2X6 U3549 ( .A(n6350), .B(n6331), .Z(n7317) );
  HS65_LL_NAND2X4 U3550 ( .A(n4282), .B(n4281), .Z(n4453) );
  HS65_LL_NAND3X5 U3551 ( .A(n7083), .B(n7082), .C(n7081), .Z(n7306) );
  HS65_LH_AOI21X2 U3552 ( .A(n8056), .B(n7697), .C(n7636), .Z(n7776) );
  HS65_LH_NOR2AX3 U3553 ( .A(n9111), .B(n7076), .Z(n7083) );
  HS65_LL_AOI21X2 U3554 ( .A(n7115), .B(n7614), .C(n7613), .Z(n8034) );
  HS65_LH_AND2X4 U3556 ( .A(\u_DataPath/jaddr_i [20]), .B(
        \u_DataPath/jaddr_i [19]), .Z(n6347) );
  HS65_LH_NOR4ABX2 U3558 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5488), .C(n5571), .D(n5353), .Z(n5372) );
  HS65_LL_OAI12X2 U3559 ( .A(n5539), .B(n5538), .C(n5537), .Z(n5593) );
  HS65_LHS_XNOR2X3 U3560 ( .A(n4045), .B(n4044), .Z(n4046) );
  HS65_LH_OAI12X3 U3561 ( .A(n3935), .B(n4929), .C(n4085), .Z(n3847) );
  HS65_LH_NOR4ABX2 U3562 ( .A(n5289), .B(n5344), .C(n5350), .D(n5288), .Z(
        n5368) );
  HS65_LH_IVX9 U3563 ( .A(\u_DataPath/jaddr_i [21]), .Z(n8163) );
  HS65_LH_IVX9 U3564 ( .A(\u_DataPath/jaddr_i [23]), .Z(n8165) );
  HS65_LH_IVX9 U3565 ( .A(write_byte), .Z(n2981) );
  HS65_LL_AOI21X2 U3566 ( .A(n4431), .B(n4363), .C(n4362), .Z(n4364) );
  HS65_LH_OAI12X3 U3568 ( .A(n4090), .B(n4929), .C(n4089), .Z(n4091) );
  HS65_LL_NOR3X4 U3569 ( .A(n5528), .B(n5527), .C(n5513), .Z(n5559) );
  HS65_LH_AOI12X2 U3573 ( .A(n5299), .B(n4017), .C(n5466), .Z(n5301) );
  HS65_LH_AOI21X2 U3574 ( .A(n5632), .B(n5630), .C(n5629), .Z(n5636) );
  HS65_LH_IVX9 U3576 ( .A(n5144), .Z(n4954) );
  HS65_LH_AOI21X2 U3577 ( .A(n5575), .B(n5015), .C(n5014), .Z(n5016) );
  HS65_LH_OAI21X2 U3578 ( .A(n5071), .B(n5070), .C(n5069), .Z(n5072) );
  HS65_LH_NAND3X5 U3579 ( .A(n5479), .B(n5478), .C(n5477), .Z(n5480) );
  HS65_LL_AOI21X2 U3580 ( .A(n5586), .B(n5009), .C(n5585), .Z(n5010) );
  HS65_LL_OAI21X2 U3583 ( .A(n5152), .B(n5616), .C(n4167), .Z(n4168) );
  HS65_LH_IVX9 U3586 ( .A(n5661), .Z(n4855) );
  HS65_LL_NOR2X6 U3589 ( .A(n4502), .B(n4863), .Z(n4951) );
  HS65_LH_AOI21X2 U3590 ( .A(n3521), .B(n4588), .C(n3830), .Z(n3831) );
  HS65_LH_IVX9 U3592 ( .A(n4939), .Z(n6123) );
  HS65_LH_AOI21X2 U3594 ( .A(n2849), .B(n4588), .C(n3904), .Z(n4496) );
  HS65_LH_AOI21X2 U3595 ( .A(n5732), .B(n5758), .C(n5731), .Z(n5799) );
  HS65_LH_IVX9 U3596 ( .A(n3935), .Z(n3482) );
  HS65_LH_AOI21X2 U3597 ( .A(n5805), .B(n5807), .C(n5734), .Z(n5735) );
  HS65_LH_IVX9 U3598 ( .A(n3426), .Z(n4502) );
  HS65_LH_NOR2X6 U3599 ( .A(n4534), .B(n4581), .Z(n5207) );
  HS65_LL_NAND2X7 U3600 ( .A(n4949), .B(n4836), .Z(n5646) );
  HS65_LH_NAND2X7 U3601 ( .A(\u_DataPath/u_idexreg/N3 ), .B(n4550), .Z(n5249)
         );
  HS65_LL_NAND2X7 U3602 ( .A(n3643), .B(n3642), .Z(n4614) );
  HS65_LL_NAND2X7 U3604 ( .A(n2851), .B(n4581), .Z(n4341) );
  HS65_LH_AOI21X2 U3605 ( .A(n6010), .B(n5936), .C(n5935), .Z(n6000) );
  HS65_LH_IVX9 U3608 ( .A(\lte_x_59/B[28] ), .Z(n4724) );
  HS65_LH_NAND2X7 U3609 ( .A(n3431), .B(n5032), .Z(n4534) );
  HS65_LL_NAND2X7 U3610 ( .A(n3490), .B(n3489), .Z(n4632) );
  HS65_LL_NOR2X6 U3611 ( .A(\lte_x_59/B[21] ), .B(n5418), .Z(n4371) );
  HS65_LH_NOR2X9 U3612 ( .A(n2840), .B(n7623), .Z(n5571) );
  HS65_LH_NAND2X7 U3613 ( .A(n5021), .B(\lte_x_59/B[16] ), .Z(n4846) );
  HS65_LH_NAND2X7 U3614 ( .A(\sub_x_53/A[20] ), .B(n4699), .Z(n4425) );
  HS65_LH_OAI12X3 U3615 ( .A(n2860), .B(n2856), .C(n3963), .Z(n4257) );
  HS65_LH_AOI21X2 U3616 ( .A(n5844), .B(n5720), .C(n5719), .Z(n5832) );
  HS65_LH_AOI21X2 U3617 ( .A(n5761), .B(n5728), .C(n5727), .Z(n5729) );
  HS65_LH_AOI21X2 U3618 ( .A(n5833), .B(n5722), .C(n5721), .Z(n5723) );
  HS65_LH_AOI21X2 U3619 ( .A(n5811), .B(n5813), .C(n5733), .Z(n5800) );
  HS65_LL_NAND2AX7 U3620 ( .A(n3546), .B(n3545), .Z(n4344) );
  HS65_LH_IVX9 U3621 ( .A(\lte_x_59/B[5] ), .Z(n5041) );
  HS65_LH_NAND2X7 U3622 ( .A(\lte_x_59/B[7] ), .B(n5030), .Z(n4624) );
  HS65_LH_IVX9 U3625 ( .A(\lte_x_59/B[26] ), .Z(n5568) );
  HS65_LL_NAND2X5 U3626 ( .A(n3474), .B(n5104), .Z(n4038) );
  HS65_LL_IVX9 U3628 ( .A(n3101), .Z(\sub_x_53/A[25] ) );
  HS65_LL_IVX18 U3632 ( .A(n3756), .Z(n4588) );
  HS65_LH_NAND2X7 U3634 ( .A(\lte_x_59/B[5] ), .B(n5040), .Z(n4107) );
  HS65_LL_NOR2AX6 U3635 ( .A(n3077), .B(n3076), .Z(\sub_x_53/A[29] ) );
  HS65_LL_NOR2X6 U3637 ( .A(\sub_x_53/A[17] ), .B(n5001), .Z(n3558) );
  HS65_LH_IVX9 U3640 ( .A(n2845), .Z(n2857) );
  HS65_LH_OAI12X3 U3642 ( .A(n8355), .B(n3409), .C(n3094), .Z(n3095) );
  HS65_LH_NOR2AX3 U3644 ( .A(n5054), .B(n2871), .Z(n4902) );
  HS65_LH_AO31X9 U3646 ( .A(n8393), .B(n2866), .C(n9376), .D(n3419), .Z(n5032)
         );
  HS65_LL_IVX4 U3648 ( .A(n4969), .Z(n3059) );
  HS65_LL_NOR2X6 U3649 ( .A(n3064), .B(n3063), .Z(\lte_x_59/B[1] ) );
  HS65_LH_NOR2X6 U3650 ( .A(n3187), .B(n3186), .Z(n3432) );
  HS65_LL_NOR2X6 U3652 ( .A(n3240), .B(n3239), .Z(n3474) );
  HS65_LL_OAI12X6 U3653 ( .A(n3192), .B(n2894), .C(n3191), .Z(n5231) );
  HS65_LL_OAI12X6 U3656 ( .A(n3224), .B(n3223), .C(n3222), .Z(n5373) );
  HS65_LL_BFX9 U3657 ( .A(n3333), .Z(n3264) );
  HS65_LH_IVX18 U3658 ( .A(n3082), .Z(n3403) );
  HS65_LL_AOI21X2 U3660 ( .A(n3404), .B(n9385), .C(n3025), .Z(n7854) );
  HS65_LH_IVX18 U3661 ( .A(n4712), .Z(n2874) );
  HS65_LLS_XOR2X3 U3665 ( .A(n2940), .B(n2846), .Z(n2964) );
  HS65_LL_NAND3X3 U3666 ( .A(n2941), .B(n7343), .C(n7089), .Z(n3052) );
  HS65_LL_IVX9 U3668 ( .A(n7084), .Z(n2846) );
  HS65_LL_NAND2X7 U3670 ( .A(\lte_x_59/B[5] ), .B(n4665), .Z(n4143) );
  HS65_LL_IVX4 U3671 ( .A(n4657), .Z(n3339) );
  HS65_LL_CBI4I1X5 U3673 ( .A(n5685), .B(n7853), .C(n7872), .D(n5684), .Z(
        n7862) );
  HS65_LL_IVX4 U3675 ( .A(n5694), .Z(n5675) );
  HS65_LL_NAND2X14 U3676 ( .A(n3308), .B(n3310), .Z(n4712) );
  HS65_LL_IVX9 U3677 ( .A(n3008), .Z(n7089) );
  HS65_LH_NAND3X2 U3680 ( .A(n7089), .B(n9031), .C(n9078), .Z(n2773) );
  HS65_LH_IVX13 U3684 ( .A(n8693), .Z(n7758) );
  HS65_LH_NAND2X2 U3685 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(nibble[0]), 
        .Z(n8575) );
  HS65_LH_IVX9 U3686 ( .A(n2988), .Z(n2801) );
  HS65_LL_NOR2AX25 U3687 ( .A(\u_DataPath/dataOut_exe_i [28]), .B(n3116), .Z(
        Address_toRAM[26]) );
  HS65_LL_NOR2AX3 U3688 ( .A(\u_DataPath/dataOut_exe_i [12]), .B(n2986), .Z(
        n3005) );
  HS65_LL_NOR2AX3 U3690 ( .A(\u_DataPath/dataOut_exe_i [10]), .B(n2986), .Z(
        n3007) );
  HS65_LH_NAND2X2 U3692 ( .A(addr_to_iram[12]), .B(addr_to_iram[13]), .Z(n7676) );
  HS65_LH_NAND2X2 U3695 ( .A(n8704), .B(addr_to_iram[15]), .Z(n7648) );
  HS65_LL_NOR2AX25 U3696 ( .A(\u_DataPath/dataOut_exe_i [13]), .B(n2986), .Z(
        Address_toRAM[11]) );
  HS65_LL_NOR2AX25 U3697 ( .A(\u_DataPath/dataOut_exe_i [27]), .B(n3116), .Z(
        Address_toRAM[25]) );
  HS65_LL_NOR2AX25 U3698 ( .A(n8728), .B(n3115), .Z(Data_in[31]) );
  HS65_LH_NOR2X2 U3702 ( .A(n5476), .B(n5522), .Z(n5515) );
  HS65_LH_OAI21X3 U3703 ( .A(n4926), .B(n3932), .C(n3934), .Z(n3477) );
  HS65_LH_CNIVX3 U3704 ( .A(n3395), .Z(n3290) );
  HS65_LH_NOR2X2 U3705 ( .A(n4724), .B(n5423), .Z(n5505) );
  HS65_LH_NAND2X2 U3706 ( .A(n2858), .B(n2864), .Z(n3871) );
  HS65_LH_CNIVX3 U3707 ( .A(n8547), .Z(n3161) );
  HS65_LH_NAND2X2 U3709 ( .A(n4717), .B(n9342), .Z(n3195) );
  HS65_LH_OAI21X3 U3710 ( .A(n4664), .B(n4637), .C(n4663), .Z(n5389) );
  HS65_LH_NOR3X1 U3711 ( .A(n5082), .B(n5081), .C(n5080), .Z(n5114) );
  HS65_LH_NAND2X2 U3715 ( .A(n4714), .B(n8518), .Z(n3254) );
  HS65_LH_NAND2X2 U3716 ( .A(\lte_x_59/B[24] ), .B(n5180), .Z(n5209) );
  HS65_LH_OAI21X3 U3717 ( .A(n5621), .B(n5620), .C(n5619), .Z(n5622) );
  HS65_LH_CNIVX3 U3719 ( .A(n3427), .Z(n5659) );
  HS65_LH_OAI21X3 U3720 ( .A(n6058), .B(n5957), .C(n5959), .Z(n5929) );
  HS65_LH_NAND2X2 U3723 ( .A(n4295), .B(n5210), .Z(n4296) );
  HS65_LH_CNIVX3 U3724 ( .A(n5405), .Z(n5476) );
  HS65_LH_IVX9 U3725 ( .A(n5618), .Z(n5241) );
  HS65_LH_NAND2X2 U3726 ( .A(\sub_x_53/A[20] ), .B(n4551), .Z(n3819) );
  HS65_LH_CNIVX3 U3727 ( .A(n5128), .Z(n3773) );
  HS65_LL_IVX2 U3728 ( .A(n4250), .Z(n5261) );
  HS65_LH_NOR2X2 U3729 ( .A(n9030), .B(n9223), .Z(n6038) );
  HS65_LH_NOR2X2 U3730 ( .A(n3905), .B(n4954), .Z(n3906) );
  HS65_LH_CNIVX3 U3731 ( .A(n5400), .Z(n5466) );
  HS65_LH_NAND2X2 U3732 ( .A(n3448), .B(n5469), .Z(n3449) );
  HS65_LH_OAI21X3 U3733 ( .A(n5627), .B(n3702), .C(n5435), .Z(n3703) );
  HS65_LH_CNIVX3 U3734 ( .A(n4230), .Z(n4303) );
  HS65_LH_AOI12X2 U3735 ( .A(\lte_x_59/B[28] ), .B(n4588), .C(n3439), .Z(n3440) );
  HS65_LH_CNIVX3 U3738 ( .A(n4849), .Z(n5203) );
  HS65_LH_NOR2X2 U3739 ( .A(n5646), .B(n5645), .Z(n5669) );
  HS65_LH_CNIVX3 U3740 ( .A(n4457), .Z(n4430) );
  HS65_LH_NAND2X2 U3742 ( .A(\u_DataPath/jaddr_i [19]), .B(n6326), .Z(n6331)
         );
  HS65_LHS_XNOR2X3 U3743 ( .A(\u_DataPath/jaddr_i [18]), .B(n8967), .Z(n7101)
         );
  HS65_LH_OAI21X3 U3744 ( .A(n5730), .B(n5759), .C(n5729), .Z(n5731) );
  HS65_LH_NAND2X2 U3745 ( .A(n7670), .B(n7649), .Z(n7650) );
  HS65_LH_CNIVX3 U3746 ( .A(n6014), .Z(n5937) );
  HS65_LH_NAND2X2 U3747 ( .A(n9185), .B(n9230), .Z(n6006) );
  HS65_LH_NAND2X2 U3748 ( .A(n9183), .B(n9232), .Z(n5978) );
  HS65_LH_NOR2X2 U3749 ( .A(n5987), .B(n5990), .Z(n5961) );
  HS65_LH_NOR2X2 U3752 ( .A(n4502), .B(n4495), .Z(n4506) );
  HS65_LH_NAND2X2 U3754 ( .A(n4084), .B(n4086), .Z(n3848) );
  HS65_LH_NOR2X2 U3755 ( .A(n7713), .B(n7711), .Z(n5168) );
  HS65_LH_NOR2X6 U3757 ( .A(n6153), .B(n6139), .Z(n6376) );
  HS65_LH_BFX9 U3758 ( .A(n9373), .Z(n7580) );
  HS65_LH_NAND3X2 U3760 ( .A(n7103), .B(n7102), .C(n7101), .Z(n7111) );
  HS65_LH_NOR2X2 U3761 ( .A(n9341), .B(n9207), .Z(n5748) );
  HS65_LH_NOR2X2 U3762 ( .A(n9181), .B(n9226), .Z(n5756) );
  HS65_LH_NAND2X2 U3763 ( .A(n9173), .B(n9231), .Z(n5876) );
  HS65_LH_CNIVX3 U3764 ( .A(n8915), .Z(n8268) );
  HS65_LH_NAND2X2 U3765 ( .A(n7659), .B(n7684), .Z(n7673) );
  HS65_LH_NOR2X2 U3766 ( .A(n7795), .B(n7794), .Z(n7307) );
  HS65_LH_NAND2X2 U3767 ( .A(n4189), .B(n8571), .Z(n4190) );
  HS65_LH_NOR2X2 U3768 ( .A(n8825), .B(n3341), .Z(n3177) );
  HS65_LH_NAND2X2 U3769 ( .A(n9173), .B(n9231), .Z(n6075) );
  HS65_LH_NAND2X2 U3770 ( .A(n8297), .B(n3407), .Z(n3104) );
  HS65_LH_NOR2X2 U3771 ( .A(n8848), .B(n3341), .Z(n3159) );
  HS65_LH_CNIVX3 U3772 ( .A(\u_DataPath/dataOut_exe_i [19]), .Z(n3188) );
  HS65_LH_OAI21X3 U3774 ( .A(n4019), .B(n3815), .C(n4018), .Z(n4020) );
  HS65_LH_OAI21X3 U3778 ( .A(n4349), .B(n4363), .C(n4949), .Z(n4095) );
  HS65_LH_NAND2X2 U3782 ( .A(n5285), .B(n4483), .Z(n4484) );
  HS65_LH_NAND2X2 U3783 ( .A(n5689), .B(n7723), .Z(n7714) );
  HS65_LH_NAND2X2 U3784 ( .A(n9039), .B(n9116), .Z(n6100) );
  HS65_LH_CNIVX3 U3785 ( .A(n7707), .Z(n7787) );
  HS65_LH_NOR2X2 U3787 ( .A(n8172), .B(\u_DataPath/immediate_ext_dec_i [4]), 
        .Z(n8076) );
  HS65_LH_NOR2X2 U3788 ( .A(n7668), .B(n7644), .Z(n7665) );
  HS65_LH_AOI12X3 U3789 ( .A(n6053), .B(n6055), .C(n5944), .Z(n5945) );
  HS65_LH_NOR2X2 U3790 ( .A(n5795), .B(n5798), .Z(n5808) );
  HS65_LH_CNIVX3 U3791 ( .A(n5799), .Z(n5868) );
  HS65_LH_NAND2X2 U3792 ( .A(n9179), .B(n9225), .Z(n5885) );
  HS65_LHS_XNOR2X3 U3793 ( .A(n9235), .B(n8268), .Z(n2980) );
  HS65_LH_NOR2X2 U3794 ( .A(n8480), .B(n7874), .Z(n7872) );
  HS65_LH_NAND2X2 U3795 ( .A(n8697), .B(n7767), .Z(n7768) );
  HS65_LH_CNIVX3 U3796 ( .A(n8235), .Z(n8287) );
  HS65_LH_CNIVX3 U3800 ( .A(n8306), .Z(n3274) );
  HS65_LHS_XNOR2X3 U3801 ( .A(n7724), .B(n7723), .Z(
        \u_DataPath/u_execute/link_value_i [14]) );
  HS65_LH_NOR2X2 U3802 ( .A(n8480), .B(n8306), .Z(n8600) );
  HS65_LH_CNIVX3 U3804 ( .A(n8394), .Z(n3412) );
  HS65_LH_NOR2X2 U3805 ( .A(n8480), .B(n8258), .Z(n8591) );
  HS65_LHS_XNOR2X3 U3806 ( .A(n7709), .B(n7708), .Z(
        \u_DataPath/u_execute/link_value_i [7]) );
  HS65_LH_MUXI21X5 U3809 ( .D0(n3175), .D1(n9383), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8385) );
  HS65_LHS_XNOR2X3 U3810 ( .A(n3517), .B(n3516), .Z(n3571) );
  HS65_LH_NOR3X1 U3811 ( .A(n7094), .B(n7093), .C(n7092), .Z(n7095) );
  HS65_LH_NAND2X2 U3812 ( .A(n9035), .B(n9115), .Z(n6049) );
  HS65_LH_CNIVX3 U3814 ( .A(n8114), .Z(n8091) );
  HS65_LH_NAND2X2 U3815 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .B(n8157), 
        .Z(n8115) );
  HS65_LH_NOR2X2 U3816 ( .A(n9082), .B(n7734), .Z(n8038) );
  HS65_LHS_XNOR2X3 U3817 ( .A(n5881), .B(n5880), .Z(\u_DataPath/toPC2_i [9])
         );
  HS65_LH_NAND2X2 U3818 ( .A(n3470), .B(\u_DataPath/cw_to_ex_i [2]), .Z(n7617)
         );
  HS65_LH_NOR2X2 U3821 ( .A(n8844), .B(n4712), .Z(n8500) );
  HS65_LH_CNIVX3 U3822 ( .A(n8600), .Z(n7974) );
  HS65_LH_AND2X4 U3823 ( .A(n3311), .B(n3310), .Z(n3312) );
  HS65_LH_CNIVX3 U3824 ( .A(n8586), .Z(n7932) );
  HS65_LH_NOR2X2 U3826 ( .A(n3062), .B(n9401), .Z(n8485) );
  HS65_LH_CNIVX3 U3827 ( .A(n8608), .Z(n8001) );
  HS65_LH_NAND3X2 U3829 ( .A(n9005), .B(n8965), .C(n8091), .Z(n8093) );
  HS65_LH_CNIVX3 U3830 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .Z(n8090) );
  HS65_LHS_XNOR2X3 U3833 ( .A(n7667), .B(n7666), .Z(\u_DataPath/pc_4_i [7]) );
  HS65_LHS_XNOR2X3 U3834 ( .A(n3125), .B(n7672), .Z(\u_DataPath/pc_4_i [15])
         );
  HS65_LH_CNIVX3 U3835 ( .A(\u_DataPath/jaddr_i [22]), .Z(n8164) );
  HS65_LH_NAND2X2 U3836 ( .A(n9084), .B(n9082), .Z(n8056) );
  HS65_LH_NAND2X2 U3837 ( .A(n7616), .B(n7615), .Z(n8160) );
  HS65_LH_OAI21X3 U3838 ( .A(n9137), .B(n8828), .C(n7847), .Z(
        \u_DataPath/dataOut_exe_i [1]) );
  HS65_LH_OAI22X1 U3840 ( .A(n9272), .B(n9270), .C(n9119), .D(n8752), .Z(
        \u_DataPath/data_read_ex_2_i [15]) );
  HS65_LH_OAI21X2 U3842 ( .A(n9189), .B(n9026), .C(n8445), .Z(
        \u_DataPath/dataOut_exe_i [29]) );
  HS65_LH_OAI22X1 U3844 ( .A(n7917), .B(n8431), .C(n7916), .D(n8430), .Z(
        \u_DataPath/data_read_ex_1_i [4]) );
  HS65_LH_OAI21X3 U3846 ( .A(n9190), .B(n8903), .C(n8312), .Z(
        \u_DataPath/dataOut_exe_i [6]) );
  HS65_LH_CNIVX3 U3848 ( .A(n8064), .Z(n8627) );
  HS65_LH_NOR2X2 U3851 ( .A(n9168), .B(n9050), .Z(\u_DataPath/u_idexreg/N16 )
         );
  HS65_LH_CNIVX3 U3853 ( .A(n8240), .Z(\u_DataPath/branch_target_i [27]) );
  HS65_LH_CNIVX3 U3854 ( .A(n8259), .Z(\u_DataPath/branch_target_i [10]) );
  HS65_LL_OR2X9 U3855 ( .A(n3411), .B(n3410), .Z(n2840) );
  HS65_LH_IVX13 U3857 ( .A(\lte_x_59/B[6] ), .Z(n2848) );
  HS65_LL_NOR2X13 U3858 ( .A(n3250), .B(n3249), .Z(n2842) );
  HS65_LL_OR2X9 U3859 ( .A(n3073), .B(n3072), .Z(n2843) );
  HS65_LL_IVX9 U3860 ( .A(\sub_x_53/A[23] ), .Z(n2860) );
  HS65_LLS_XNOR2X3 U3861 ( .A(n4160), .B(n4159), .Z(n2844) );
  HS65_LL_AND2X18 U3862 ( .A(n5136), .B(n3401), .Z(n2845) );
  HS65_LL_NOR3X4 U3864 ( .A(n5165), .B(n5164), .C(n5683), .Z(n7852) );
  HS65_LL_NAND3AX13 U3865 ( .A(n2939), .B(n2938), .C(n2937), .Z(n3308) );
  HS65_LL_NAND2X4 U3867 ( .A(n8468), .B(n8465), .Z(n4790) );
  HS65_LL_AOI12X6 U3868 ( .A(n7631), .B(n4174), .C(n4173), .Z(n8465) );
  HS65_LL_NAND3X3 U3869 ( .A(n4857), .B(n4744), .C(n4743), .Z(n4745) );
  HS65_LL_NAND3X5 U3871 ( .A(n5561), .B(n5560), .C(n5559), .Z(n5591) );
  HS65_LL_AOI12X2 U3874 ( .A(n5606), .B(n3499), .C(n3498), .Z(n3500) );
  HS65_LL_NOR2X6 U3878 ( .A(n3320), .B(n3319), .Z(\lte_x_59/B[6] ) );
  HS65_LL_NAND2X5 U3879 ( .A(n4365), .B(n4364), .Z(n4366) );
  HS65_LL_NAND3X5 U3880 ( .A(n4361), .B(n4360), .C(n4359), .Z(n4362) );
  HS65_LL_NAND2AX7 U3881 ( .A(n3551), .B(n2899), .Z(n4886) );
  HS65_LL_NOR2X3 U3882 ( .A(n4755), .B(n4754), .Z(n4756) );
  HS65_LL_NAND3X5 U3883 ( .A(n3487), .B(n3486), .C(n4593), .Z(n3490) );
  HS65_LL_BFX9 U3885 ( .A(n3432), .Z(n2849) );
  HS65_LL_OAI12X2 U3886 ( .A(n3366), .B(n5179), .C(n4940), .Z(n4941) );
  HS65_LH_OAI112X3 U3887 ( .A(n5334), .B(n5301), .C(n5405), .D(n5479), .Z(
        n5308) );
  HS65_LL_NOR2X6 U3888 ( .A(\lte_x_59/B[1] ), .B(n4805), .Z(n4823) );
  HS65_LLS_XNOR2X3 U3889 ( .A(\lte_x_59/B[1] ), .B(n4805), .Z(n4808) );
  HS65_LL_IVX9 U3890 ( .A(n2840), .Z(n2851) );
  HS65_LL_NOR2X3 U3891 ( .A(n8355), .B(n9401), .Z(n8525) );
  HS65_LL_NOR2X3 U3892 ( .A(n5241), .B(n5240), .Z(n5242) );
  HS65_LL_NOR2X6 U3896 ( .A(n3770), .B(n3769), .Z(n4522) );
  HS65_LL_AOI12X2 U3897 ( .A(n4587), .B(\lte_x_59/B[15] ), .C(n3982), .Z(n3983) );
  HS65_LL_NAND2X5 U3898 ( .A(\lte_x_59/B[4] ), .B(n5032), .Z(n4477) );
  HS65_LL_OAI21X3 U3899 ( .A(n5646), .B(n4180), .C(n3660), .Z(n3661) );
  HS65_LL_OAI211X3 U3900 ( .A(n5226), .B(n5646), .C(n4586), .D(n4585), .Z(
        n4602) );
  HS65_LL_NOR2X6 U3901 ( .A(n3773), .B(n3772), .Z(n4513) );
  HS65_LL_AOI12X2 U3902 ( .A(n5526), .B(n5525), .C(n5524), .Z(n5538) );
  HS65_LL_OAI21X3 U3903 ( .A(n5485), .B(n5337), .C(n5336), .Z(n5338) );
  HS65_LL_AOI12X2 U3906 ( .A(n4551), .B(n3521), .C(n4153), .Z(n3455) );
  HS65_LL_IVX9 U3907 ( .A(n3521), .Z(n4671) );
  HS65_LL_IVX9 U3908 ( .A(n4966), .Z(n2873) );
  HS65_LL_NAND2X14 U3909 ( .A(n3967), .B(n2872), .Z(n5152) );
  HS65_LL_IVX9 U3912 ( .A(\sub_x_53/A[20] ), .Z(n4700) );
  HS65_LLS_XNOR2X3 U3913 ( .A(\sub_x_53/A[20] ), .B(n4699), .Z(n4768) );
  HS65_LL_AOI12X2 U3915 ( .A(\lte_x_59/B[7] ), .B(n4588), .C(n3670), .Z(n3920)
         );
  HS65_LL_IVX2 U3916 ( .A(\lte_x_59/B[7] ), .Z(n5031) );
  HS65_LL_NOR2X13 U3917 ( .A(n3200), .B(n3199), .Z(\sub_x_53/A[17] ) );
  HS65_LH_IVX13 U3918 ( .A(n5568), .Z(n2853) );
  HS65_LL_IVX9 U3919 ( .A(\lte_x_59/B[26] ), .Z(n2854) );
  HS65_LL_NAND2X7 U3920 ( .A(n4970), .B(n4974), .Z(n5423) );
  HS65_LL_OAI211X1 U3921 ( .A(n5572), .B(n5571), .C(n5570), .D(n5569), .Z(
        n5573) );
  HS65_LL_NOR2X3 U3922 ( .A(n5571), .B(n4230), .Z(n5453) );
  HS65_LL_OAI21X2 U3923 ( .A(n5450), .B(n5571), .C(n5449), .Z(n5451) );
  HS65_LL_AOI112X4 U3925 ( .A(\lte_x_59/B[21] ), .B(n4351), .C(n3667), .D(
        n3666), .Z(n4185) );
  HS65_LL_AOI12X2 U3926 ( .A(\lte_x_59/B[21] ), .B(n4544), .C(n3903), .Z(n4497) );
  HS65_LL_OAI21X2 U3928 ( .A(n5388), .B(n5387), .C(n4143), .Z(n5391) );
  HS65_LL_IVX9 U3932 ( .A(n2843), .Z(n2858) );
  HS65_LL_IVX9 U3933 ( .A(n4674), .Z(n5376) );
  HS65_LL_NAND3X5 U3934 ( .A(n3837), .B(n3836), .C(n3835), .Z(n4839) );
  HS65_LL_AOI12X6 U3935 ( .A(n3618), .B(n4879), .C(n3617), .Z(n5610) );
  HS65_LLS_XNOR2X3 U3936 ( .A(n2849), .B(n5231), .Z(n5232) );
  HS65_LLS_XNOR2X3 U3937 ( .A(\sub_x_53/A[0] ), .B(n5136), .Z(n5141) );
  HS65_LL_IVX4 U3941 ( .A(n5691), .Z(n3224) );
  HS65_LL_OAI21X2 U3942 ( .A(n4573), .B(n5383), .C(n5090), .Z(n5384) );
  HS65_LL_AOI12X6 U3943 ( .A(n5672), .B(n5671), .C(n5670), .Z(n5673) );
  HS65_LL_AOI12X2 U3945 ( .A(\lte_x_59/B[4] ), .B(n4551), .C(n3400), .Z(n3875)
         );
  HS65_LLS_XNOR2X3 U3947 ( .A(\lte_x_59/B[8] ), .B(n5373), .Z(n4762) );
  HS65_LL_NOR2X6 U3949 ( .A(\lte_x_59/B[5] ), .B(n5040), .Z(n4105) );
  HS65_LL_NAND2X4 U3950 ( .A(\lte_x_59/B[5] ), .B(n2864), .Z(n4542) );
  HS65_LL_NAND2X5 U3951 ( .A(n3379), .B(n5632), .Z(n3375) );
  HS65_LL_NAND2X7 U3952 ( .A(n3751), .B(n3383), .Z(n4330) );
  HS65_LL_OAI21X3 U3953 ( .A(n5405), .B(n4049), .C(n4050), .Z(n4917) );
  HS65_LL_IVX4 U3954 ( .A(n3474), .Z(n5105) );
  HS65_LL_NAND2X4 U3957 ( .A(n4385), .B(n4382), .Z(n4121) );
  HS65_LL_NAND2X4 U3959 ( .A(n4836), .B(n4886), .Z(n4382) );
  HS65_LL_AOI12X2 U3960 ( .A(\lte_x_59/B[6] ), .B(n4588), .C(n3764), .Z(n3765)
         );
  HS65_LL_NAND3X3 U3963 ( .A(n8429), .B(n8875), .C(n8896), .Z(
        \u_DataPath/dataOut_exe_i [0]) );
  HS65_LH_NAND2X2 U3964 ( .A(\u_DataPath/u_execute/ovf_i ), .B(n2733), .Z(
        n8423) );
  HS65_LL_OAI12X3 U3967 ( .A(n9189), .B(n8901), .C(n8416), .Z(
        \u_DataPath/dataOut_exe_i [28]) );
  HS65_LL_OAI12X3 U3969 ( .A(n9190), .B(n8900), .C(n8328), .Z(
        \u_DataPath/dataOut_exe_i [25]) );
  HS65_LL_NAND2X4 U3970 ( .A(n8419), .B(n8899), .Z(
        \u_DataPath/dataOut_exe_i [31]) );
  HS65_LL_OAI12X3 U3971 ( .A(n9189), .B(n8891), .C(n8359), .Z(
        \u_DataPath/dataOut_exe_i [23]) );
  HS65_LL_CNIVX3 U3972 ( .A(n5598), .Z(n5599) );
  HS65_LL_AOI12X4 U3973 ( .A(n5285), .B(n3628), .C(n3627), .Z(n8478) );
  HS65_LL_OAI12X3 U3974 ( .A(n5602), .B(n5598), .C(n4243), .Z(n7841) );
  HS65_LL_NAND3X2 U3975 ( .A(n3569), .B(n3568), .C(n3567), .Z(n3570) );
  HS65_LL_IVX2 U3977 ( .A(n8464), .Z(n4793) );
  HS65_LH_NAND2AX7 U3980 ( .A(n5705), .B(n5704), .Z(n5706) );
  HS65_LL_OAI21X2 U3983 ( .A(n5633), .B(n3636), .C(n3635), .Z(n3637) );
  HS65_LL_OAI21X2 U3984 ( .A(n3806), .B(n2859), .C(n3805), .Z(n3807) );
  HS65_LH_NOR2X6 U3985 ( .A(n5490), .B(n5489), .Z(n5494) );
  HS65_LH_IVX4 U3986 ( .A(n2859), .Z(n4297) );
  HS65_LH_AOI21X6 U3987 ( .A(n5195), .B(n4238), .C(n4237), .Z(n4239) );
  HS65_LH_NOR2X5 U3988 ( .A(n4995), .B(n4994), .Z(n5118) );
  HS65_LH_IVX4 U3990 ( .A(n4948), .Z(n4533) );
  HS65_LH_CNIVX3 U3991 ( .A(n5250), .Z(n5251) );
  HS65_LH_AOI12X2 U3992 ( .A(n3389), .B(n5195), .C(n3388), .Z(n3390) );
  HS65_LH_IVX7 U3993 ( .A(n4236), .Z(n4237) );
  HS65_LH_NAND2X2 U3994 ( .A(n4512), .B(n5614), .Z(n4150) );
  HS65_LL_NAND2X2 U3995 ( .A(n5615), .B(n4388), .Z(n4405) );
  HS65_LH_IVX7 U3996 ( .A(n5616), .Z(n5623) );
  HS65_LH_AOI21X4 U3997 ( .A(n5029), .B(n5020), .C(n5019), .Z(n5078) );
  HS65_LH_IVX18 U3998 ( .A(n4879), .Z(n4929) );
  HS65_LH_AOI31X3 U3999 ( .A(n5582), .B(n5581), .C(n5580), .D(n5579), .Z(n5589) );
  HS65_LH_NAND3X5 U4001 ( .A(n4431), .B(n5321), .C(n4430), .Z(n3469) );
  HS65_LL_NAND3X3 U4003 ( .A(n4010), .B(n4009), .C(n4008), .Z(n4536) );
  HS65_LH_CNIVX3 U4004 ( .A(n4816), .Z(n4830) );
  HS65_LH_NAND2X7 U4005 ( .A(n5208), .B(n5210), .Z(n3621) );
  HS65_LH_AOI13X3 U4006 ( .A(n4845), .B(n4879), .C(n3618), .D(n3561), .Z(n3562) );
  HS65_LH_NOR2X3 U4007 ( .A(n5201), .B(n5200), .Z(n5202) );
  HS65_LH_NAND2X4 U4008 ( .A(n4086), .B(n3482), .Z(n4090) );
  HS65_LH_AOI12X2 U4009 ( .A(n5309), .B(n5308), .C(n5307), .Z(n5339) );
  HS65_LH_OAI12X3 U4010 ( .A(n5646), .B(n3966), .C(n3965), .Z(n3977) );
  HS65_LH_IVX4 U4012 ( .A(n4606), .Z(n3727) );
  HS65_LH_IVX4 U4014 ( .A(n5194), .Z(n5197) );
  HS65_LH_NAND2X7 U4015 ( .A(n5192), .B(n5194), .Z(n3578) );
  HS65_LH_NAND2X5 U4016 ( .A(n3426), .B(n4164), .Z(n5616) );
  HS65_LH_NAND2X7 U4017 ( .A(n4930), .B(n3482), .Z(n4931) );
  HS65_LH_OAI21X3 U4018 ( .A(n5226), .B(n3427), .C(n3711), .Z(n3730) );
  HS65_LH_NOR2X6 U4019 ( .A(n5528), .B(n5527), .Z(n5584) );
  HS65_LH_NOR2X6 U4020 ( .A(n3606), .B(n3605), .Z(n3607) );
  HS65_LH_NAND2X5 U4021 ( .A(n3389), .B(n5194), .Z(n3391) );
  HS65_LH_NAND2X5 U4022 ( .A(n4270), .B(n4269), .Z(n4271) );
  HS65_LH_OAI12X3 U4024 ( .A(n4855), .B(n5620), .C(n4268), .Z(n4274) );
  HS65_LH_OAI12X3 U4025 ( .A(n4855), .B(n4522), .C(n4521), .Z(n4532) );
  HS65_LH_AOI21X2 U4026 ( .A(n4942), .B(n4839), .C(n3857), .Z(n3886) );
  HS65_LH_OAI21X3 U4027 ( .A(n4803), .B(n5176), .C(n4133), .Z(n4137) );
  HS65_LH_NOR2X5 U4028 ( .A(n4232), .B(n4330), .Z(n4238) );
  HS65_LH_NAND2X5 U4029 ( .A(n5306), .B(n5305), .Z(n5307) );
  HS65_LH_NAND2X7 U4030 ( .A(n5520), .B(n5515), .Z(n5541) );
  HS65_LH_NOR2X6 U4031 ( .A(n5146), .B(n3858), .Z(n3859) );
  HS65_LH_OAI21X3 U4032 ( .A(n5177), .B(n4838), .C(n4837), .Z(n4844) );
  HS65_LH_NOR2X5 U4033 ( .A(n5018), .B(n5000), .Z(n5029) );
  HS65_LH_NAND3X5 U4034 ( .A(n3776), .B(n3775), .C(n3774), .Z(n3777) );
  HS65_LH_NAND2X5 U4035 ( .A(n5659), .B(n5206), .Z(n3428) );
  HS65_LH_NOR2X2 U4037 ( .A(n4673), .B(n4684), .Z(n4694) );
  HS65_LH_OAI21X3 U4038 ( .A(n4730), .B(n4729), .C(n4728), .Z(n4731) );
  HS65_LH_IVX4 U4040 ( .A(n5542), .Z(n5106) );
  HS65_LH_IVX9 U4041 ( .A(n4330), .Z(n3389) );
  HS65_LH_NAND2X4 U4043 ( .A(n5564), .B(n5346), .Z(n5350) );
  HS65_LH_NAND2X5 U4044 ( .A(n4497), .B(n4496), .Z(n4616) );
  HS65_LH_NAND2X4 U4045 ( .A(n3426), .B(n4344), .Z(n3587) );
  HS65_LL_CNIVX3 U4046 ( .A(n5211), .Z(n5212) );
  HS65_LH_AO12X9 U4048 ( .A(n4041), .B(n4040), .C(n4039), .Z(n4042) );
  HS65_LH_IVX9 U4050 ( .A(n4515), .Z(n5620) );
  HS65_LH_IVX4 U4051 ( .A(n4610), .Z(n3865) );
  HS65_LH_NOR2X5 U4052 ( .A(n4954), .B(n3555), .Z(n4874) );
  HS65_LH_NAND3X3 U4054 ( .A(n3426), .B(n5672), .C(n4344), .Z(n3581) );
  HS65_LH_NOR2X5 U4055 ( .A(n5241), .B(n5172), .Z(n3438) );
  HS65_LH_IVX4 U4057 ( .A(n4304), .Z(n4307) );
  HS65_LHS_XOR2X6 U4058 ( .A(n4574), .B(n4540), .Z(n4569) );
  HS65_LH_NAND3X5 U4059 ( .A(n2864), .B(n6123), .C(n4806), .Z(n4807) );
  HS65_LH_OAI21X3 U4060 ( .A(n5176), .B(n5135), .C(n5134), .Z(n5150) );
  HS65_LH_NAND2X4 U4061 ( .A(n5618), .B(n5644), .Z(n4521) );
  HS65_LH_IVX7 U4062 ( .A(n5644), .Z(n5645) );
  HS65_LH_NAND2X7 U4063 ( .A(n4211), .B(n4290), .Z(n4220) );
  HS65_LH_IVX4 U4064 ( .A(n4497), .Z(n4498) );
  HS65_LH_CNIVX3 U4065 ( .A(n4500), .Z(n4501) );
  HS65_LH_NOR2X6 U4066 ( .A(n4924), .B(n3936), .Z(n3939) );
  HS65_LH_IVX9 U4067 ( .A(n5274), .Z(n4245) );
  HS65_LH_IVX7 U4068 ( .A(n4016), .Z(n3950) );
  HS65_LH_NOR3X2 U4070 ( .A(n4502), .B(n5152), .C(n4197), .Z(n4028) );
  HS65_LH_NAND2X5 U4071 ( .A(n5270), .B(n3197), .Z(n5279) );
  HS65_LH_NOR3X4 U4072 ( .A(n3783), .B(n3820), .C(n3782), .Z(n4526) );
  HS65_LH_IVX4 U4075 ( .A(n4702), .Z(n4703) );
  HS65_LH_NAND2X5 U4076 ( .A(n5286), .B(n5572), .Z(n5287) );
  HS65_LH_NAND2X7 U4077 ( .A(n5572), .B(n4727), .Z(n4730) );
  HS65_LH_IVX7 U4078 ( .A(n5507), .Z(n5510) );
  HS65_LH_IVX4 U4079 ( .A(n4761), .Z(n3451) );
  HS65_LH_NOR2X3 U4081 ( .A(n4939), .B(n4938), .Z(n4946) );
  HS65_LH_NOR2X2 U4082 ( .A(n5421), .B(n5441), .Z(n5429) );
  HS65_LH_OAI31X5 U4083 ( .A(n5133), .B(n5139), .C(n5132), .D(n5131), .Z(n5134) );
  HS65_LH_IVX7 U4085 ( .A(n4488), .Z(n4489) );
  HS65_LH_AOI21X6 U4086 ( .A(\lte_x_59/B[28] ), .B(n2864), .C(n3548), .Z(n3586) );
  HS65_LH_IVX4 U4088 ( .A(n4930), .Z(n3936) );
  HS65_LH_IVX7 U4089 ( .A(n5269), .Z(n3197) );
  HS65_LH_NAND2X4 U4091 ( .A(n3559), .B(n3472), .Z(n3565) );
  HS65_LH_NOR2X6 U4092 ( .A(\lte_x_59/B[28] ), .B(n5423), .Z(n4320) );
  HS65_LH_NOR2X2 U4093 ( .A(n4630), .B(n4626), .Z(n4633) );
  HS65_LH_NAND2X4 U4094 ( .A(n3474), .B(n2864), .Z(n4590) );
  HS65_LH_NAND2X7 U4095 ( .A(n4930), .B(n3478), .Z(n3481) );
  HS65_LH_AOI21X4 U4096 ( .A(n3478), .B(n4927), .C(n3477), .Z(n3479) );
  HS65_LH_NOR2X6 U4097 ( .A(n3474), .B(n3359), .Z(n3949) );
  HS65_LH_IVX7 U4098 ( .A(n3819), .Z(n3824) );
  HS65_LH_NAND2X5 U4100 ( .A(n3832), .B(n3956), .Z(n3460) );
  HS65_LH_OAI12X3 U4101 ( .A(n5356), .B(n5363), .C(n5292), .Z(n5586) );
  HS65_LH_NAND2X7 U4102 ( .A(n3763), .B(n5127), .Z(n3766) );
  HS65_LH_IVX4 U4104 ( .A(n3840), .Z(n3768) );
  HS65_LH_NAND2X4 U4106 ( .A(n5234), .B(n5233), .Z(n5235) );
  HS65_LH_NAND2X5 U4107 ( .A(n5256), .B(n5255), .Z(n5265) );
  HS65_LH_OAI12X3 U4108 ( .A(n3749), .B(n3629), .C(n5443), .Z(n5444) );
  HS65_LH_NAND2X2 U4109 ( .A(n4373), .B(n4372), .Z(n4379) );
  HS65_LH_IVX9 U4110 ( .A(n5319), .Z(n5465) );
  HS65_LH_NOR2X5 U4112 ( .A(n4765), .B(n4764), .Z(n4766) );
  HS65_LH_NAND2X7 U4113 ( .A(\lte_x_59/B[28] ), .B(n3129), .Z(n4331) );
  HS65_LH_IVX4 U4116 ( .A(n3838), .Z(n3434) );
  HS65_LH_NOR2X5 U4117 ( .A(n4742), .B(n4741), .Z(n4743) );
  HS65_LH_OAI21X3 U4120 ( .A(n4795), .B(n4671), .C(n4062), .Z(n3645) );
  HS65_LH_IVX9 U4121 ( .A(n4507), .Z(n4197) );
  HS65_LH_OAI12X3 U4123 ( .A(n4675), .B(n5129), .C(n3644), .Z(n3646) );
  HS65_LH_NOR2X5 U4125 ( .A(n4682), .B(n5129), .Z(n4156) );
  HS65_LH_IVX4 U4126 ( .A(n4034), .Z(n4035) );
  HS65_LH_NAND2X7 U4127 ( .A(\lte_x_59/B[9] ), .B(n4587), .Z(n3870) );
  HS65_LH_NAND2X5 U4128 ( .A(\lte_x_59/B[22] ), .B(n4551), .Z(n3963) );
  HS65_LH_CNIVX3 U4130 ( .A(n5254), .Z(n5255) );
  HS65_LH_IVX4 U4131 ( .A(n5232), .Z(n5233) );
  HS65_LH_IVX4 U4132 ( .A(n4084), .Z(n4088) );
  HS65_LH_CNIVX3 U4133 ( .A(n4371), .Z(n4372) );
  HS65_LH_NAND2X5 U4134 ( .A(\sub_x_53/A[30] ), .B(n4966), .Z(n4289) );
  HS65_LH_NAND2AX7 U4136 ( .A(n5320), .B(n2864), .Z(n5127) );
  HS65_LL_OAI21X2 U4137 ( .A(n5258), .B(n5254), .C(n5256), .Z(n3496) );
  HS65_LH_NAND2X4 U4138 ( .A(\lte_x_59/B[4] ), .B(n4544), .Z(n3763) );
  HS65_LH_IVX4 U4139 ( .A(n4924), .Z(n4925) );
  HS65_LH_IVX4 U4142 ( .A(n3800), .Z(n3801) );
  HS65_LH_NOR2X6 U4143 ( .A(n4711), .B(n5129), .Z(n3548) );
  HS65_LH_IVX4 U4144 ( .A(n5509), .Z(n5364) );
  HS65_LH_NAND2X7 U4145 ( .A(\sub_x_53/A[30] ), .B(n4587), .Z(n3544) );
  HS65_LH_NOR2X6 U4146 ( .A(n4637), .B(n4643), .Z(n3353) );
  HS65_LH_NOR2X5 U4147 ( .A(n4700), .B(n4699), .Z(n5471) );
  HS65_LH_NOR2X3 U4148 ( .A(n4986), .B(n5005), .Z(n5355) );
  HS65_LH_IVX9 U4149 ( .A(n5531), .Z(n5511) );
  HS65_LH_IVX4 U4150 ( .A(n4740), .Z(n4741) );
  HS65_LH_NAND2X4 U4153 ( .A(n5004), .B(n5231), .Z(n5534) );
  HS65_LH_IVX9 U4154 ( .A(n4672), .Z(n5294) );
  HS65_LH_IVX7 U4155 ( .A(n5396), .Z(n5335) );
  HS65_LH_NAND2X5 U4156 ( .A(n4671), .B(n5048), .Z(n5516) );
  HS65_LH_IVX4 U4158 ( .A(n4768), .Z(n4441) );
  HS65_LH_NAND2X4 U4159 ( .A(\lte_x_59/B[16] ), .B(n4551), .Z(n3839) );
  HS65_LH_NOR2X3 U4161 ( .A(n3529), .B(n5022), .Z(n4850) );
  HS65_LH_IVX9 U4162 ( .A(n5193), .Z(n3576) );
  HS65_LH_IVX7 U4163 ( .A(n4774), .Z(n3610) );
  HS65_LH_NAND2X5 U4164 ( .A(n5397), .B(n3231), .Z(n3853) );
  HS65_LH_NAND2X5 U4165 ( .A(\lte_x_59/B[16] ), .B(n4985), .Z(n5506) );
  HS65_LH_NAND2X7 U4166 ( .A(\u_DataPath/u_idexreg/N3 ), .B(n4512), .Z(n4939)
         );
  HS65_LH_IVX18 U4168 ( .A(n4726), .Z(\sub_x_53/A[30] ) );
  HS65_LL_NOR2X2 U4169 ( .A(\lte_x_59/B[24] ), .B(n3382), .Z(n3575) );
  HS65_LH_NAND2AX7 U4170 ( .A(\lte_x_59/B[14] ), .B(n5061), .Z(n4672) );
  HS65_LH_IVX4 U4172 ( .A(n5095), .Z(n5096) );
  HS65_LH_IVX4 U4173 ( .A(n5327), .Z(n5097) );
  HS65_LL_BFX9 U4175 ( .A(n3547), .Z(\sub_x_53/A[27] ) );
  HS65_LH_NAND2X7 U4176 ( .A(n2853), .B(n3384), .Z(n3749) );
  HS65_LH_IVX4 U4177 ( .A(n4573), .Z(n4661) );
  HS65_LL_NAND2X4 U4179 ( .A(\lte_x_59/B[18] ), .B(n5005), .Z(n5258) );
  HS65_LH_NOR2X5 U4180 ( .A(n2849), .B(n5231), .Z(n5254) );
  HS65_LH_NAND2X4 U4181 ( .A(n4624), .B(n4623), .Z(n4635) );
  HS65_LL_CNBFX10 U4182 ( .A(n2856), .Z(n4583) );
  HS65_LL_IVX18 U4184 ( .A(n3756), .Z(n4551) );
  HS65_LH_OAI22X4 U4185 ( .A(n7096), .B(n8353), .C(n7900), .D(n8349), .Z(
        \u_DataPath/data_read_ex_2_i [22]) );
  HS65_LH_OAI22X4 U4186 ( .A(n7096), .B(n8343), .C(n7900), .D(n8338), .Z(
        \u_DataPath/data_read_ex_2_i [13]) );
  HS65_LH_OAI22X4 U4187 ( .A(n7096), .B(n8348), .C(n7900), .D(n8344), .Z(
        \u_DataPath/data_read_ex_2_i [11]) );
  HS65_LH_OAI22X4 U4188 ( .A(n7096), .B(n8337), .C(n7900), .D(n8331), .Z(
        \u_DataPath/data_read_ex_2_i [9]) );
  HS65_LL_NOR2X6 U4190 ( .A(n3061), .B(n3060), .Z(\lte_x_59/B[21] ) );
  HS65_LH_IVX7 U4191 ( .A(n4769), .Z(n4553) );
  HS65_LL_NOR2X6 U4194 ( .A(n3266), .B(n3265), .Z(n3521) );
  HS65_LH_CNIVX3 U4195 ( .A(n4596), .Z(n4561) );
  HS65_LL_IVX4 U4196 ( .A(n5104), .Z(n3359) );
  HS65_LH_IVX18 U4199 ( .A(n5652), .Z(\lte_x_59/B[22] ) );
  HS65_LH_IVX18 U4200 ( .A(n5054), .Z(\lte_x_59/B[9] ) );
  HS65_LH_OAI22X6 U4201 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [27]), .C(
        n8374), .D(n3409), .Z(n3107) );
  HS65_LH_NOR2X3 U4204 ( .A(n9167), .B(n8916), .Z(\u_DataPath/cw_exmem_i [4])
         );
  HS65_LL_NOR2X3 U4205 ( .A(n3118), .B(n7770), .Z(n7780) );
  HS65_LL_NAND3X5 U4206 ( .A(n2903), .B(n3081), .C(n3080), .Z(n5054) );
  HS65_LHS_XOR2X3 U4207 ( .A(n3118), .B(n7770), .Z(\u_DataPath/pc_4_i [28]) );
  HS65_LL_NAND2X5 U4209 ( .A(n8272), .B(n8298), .Z(n8452) );
  HS65_LH_AO22X9 U4210 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ), .D(
        n7586), .Z(n6335) );
  HS65_LH_AO22X9 U4211 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ), .D(
        n7318), .Z(n6336) );
  HS65_LH_AO22X9 U4212 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ), .B(n7578), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ), .Z(n7037)
         );
  HS65_LH_AO22X9 U4214 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ), .D(
        n7318), .Z(n7041) );
  HS65_LH_AO22X9 U4215 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ), .B(n7578), 
        .C(n7310), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ), .Z(n7017) );
  HS65_LH_AOI22X3 U4216 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ), .D(
        n6625), .Z(n7129) );
  HS65_LH_AOI22X3 U4219 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ), .D(
        n6624), .Z(n7130) );
  HS65_LH_AOI22X3 U4220 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ), .B(n7525), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ), .Z(n6343)
         );
  HS65_LH_AO22X9 U4222 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ), .D(n7318), .Z(n7021) );
  HS65_LH_AO22X9 U4223 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ), .D(
        n7318), .Z(n6749) );
  HS65_LH_AOI22X3 U4224 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ), .D(
        n2891), .Z(n6674) );
  HS65_LH_AOI22X3 U4226 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ), .Z(n7606)
         );
  HS65_LH_AO22X9 U4227 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ), .D(
        n7318), .Z(n7322) );
  HS65_LH_AOI22X3 U4228 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ), .D(
        n6625), .Z(n6231) );
  HS65_LH_AOI22X3 U4229 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ), .Z(n7531)
         );
  HS65_LH_AO22X9 U4230 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ), .D(
        n7318), .Z(n7209) );
  HS65_LH_AOI22X3 U4234 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ), .D(n6957), .Z(n6705) );
  HS65_LH_AOI22X3 U4237 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ), .D(
        n6957), .Z(n6678) );
  HS65_LH_AO22X9 U4238 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ), .D(n7318), .Z(n6772) );
  HS65_LH_AOI22X3 U4239 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ), .D(n6957), .Z(n6773) );
  HS65_LH_AOI22X3 U4240 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ), .D(
        n6957), .Z(n6813) );
  HS65_LH_AOI22X3 U4241 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ), .Z(n7551)
         );
  HS65_LH_AOI22X3 U4242 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ), .Z(n7485)
         );
  HS65_LH_AOI22X3 U4245 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ), .Z(n6962)
         );
  HS65_LH_AO22X9 U4246 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ), .D(
        n7318), .Z(n7189) );
  HS65_LH_AOI22X3 U4247 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ), .Z(n7571)
         );
  HS65_LH_AO22X9 U4249 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ), .B(n7578), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ), .Z(n7057)
         );
  HS65_LH_AO22X9 U4251 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ), .D(
        n7318), .Z(n7061) );
  HS65_LH_AOI22X3 U4253 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ), .D(
        n7285), .Z(n6639) );
  HS65_LH_AO22X9 U4254 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ), .D(
        n7282), .Z(n6641) );
  HS65_LH_AOI22X3 U4255 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ), .Z(n7465)
         );
  HS65_LH_AO22X9 U4257 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ), .D(
        n7318), .Z(n7001) );
  HS65_LH_AO22X9 U4258 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ), .B(n7578), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ), .Z(n6997)
         );
  HS65_LH_AOI22X3 U4262 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ), .D(
        n6957), .Z(n6793) );
  HS65_LH_AOI22X3 U4263 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ), .D(n6957), .Z(n6725) );
  HS65_LH_AOI22X3 U4265 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ), .D(
        n6625), .Z(n6136) );
  HS65_LH_AO22X9 U4267 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ), .D(
        n7318), .Z(n6792) );
  HS65_LH_AO22X9 U4268 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ), .D(
        n7318), .Z(n6981) );
  HS65_LH_AOI22X4 U4272 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ), .Z(n7409)
         );
  HS65_LH_AOI22X4 U4273 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][30] ), .Z(n7410)
         );
  HS65_LH_AO22X9 U4275 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ), .D(n7318), .Z(n6724) );
  HS65_LH_AOI22X3 U4276 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ), .Z(n7445)
         );
  HS65_LH_AOI22X3 U4277 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ), .D(
        n2891), .Z(n6722) );
  HS65_LH_AO22X9 U4278 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ), .D(n7318), .Z(n7249) );
  HS65_LH_AO22X9 U4279 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ), .D(
        n6629), .Z(n7166) );
  HS65_LL_AOI12X4 U4280 ( .A(n6105), .B(n6107), .C(n5941), .Z(n5974) );
  HS65_LL_OAI12X2 U4282 ( .A(n8266), .B(n3340), .C(n3104), .Z(n3105) );
  HS65_LH_IVX9 U4283 ( .A(n8497), .Z(n3323) );
  HS65_LH_NOR2X6 U4284 ( .A(n8867), .B(n3341), .Z(n3342) );
  HS65_LH_NOR2X6 U4285 ( .A(n3275), .B(n8522), .Z(n3276) );
  HS65_LH_NOR2X2 U4286 ( .A(rst), .B(n8554), .Z(
        \u_DataPath/mem_writedata_out_i [25]) );
  HS65_LH_NOR2X6 U4289 ( .A(n8861), .B(n3341), .Z(n3064) );
  HS65_LL_NAND3X3 U4291 ( .A(n8135), .B(n8134), .C(n8318), .Z(n8301) );
  HS65_LL_IVX9 U4293 ( .A(n4712), .Z(n3291) );
  HS65_LH_NOR2X6 U4294 ( .A(n3274), .B(n7868), .Z(n8522) );
  HS65_LH_NAND2X5 U4295 ( .A(n4714), .B(n8524), .Z(n3275) );
  HS65_LH_NOR2X6 U4296 ( .A(n8243), .B(n7868), .Z(n8547) );
  HS65_LH_NAND2X4 U4297 ( .A(n8044), .B(n8043), .Z(opcode_i[0]) );
  HS65_LH_NAND2X5 U4298 ( .A(n4714), .B(n8553), .Z(n3141) );
  HS65_LH_NAND2X4 U4299 ( .A(n8044), .B(n8036), .Z(opcode_i[2]) );
  HS65_LL_NOR2X3 U4302 ( .A(n3119), .B(n7759), .Z(n7704) );
  HS65_LH_BFX18 U4303 ( .A(n8483), .Z(n7922) );
  HS65_LL_AOI12X4 U4305 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n8573), .C(
        n8133), .Z(n8318) );
  HS65_LH_BFX18 U4306 ( .A(n8483), .Z(n7923) );
  HS65_LH_AOI21X6 U4308 ( .A(n2896), .B(n3299), .C(n3298), .Z(n3300) );
  HS65_LH_NAND2X7 U4309 ( .A(n3260), .B(n2866), .Z(n8514) );
  HS65_LH_NAND2X7 U4310 ( .A(n2896), .B(n3257), .Z(n6125) );
  HS65_LH_NAND2X4 U4312 ( .A(n3307), .B(n3407), .Z(n3304) );
  HS65_LH_NOR2X5 U4313 ( .A(n7854), .B(n9401), .Z(n8528) );
  HS65_LH_NOR2X6 U4315 ( .A(\u_DataPath/dataOut_exe_i [21]), .B(n8390), .Z(
        n8541) );
  HS65_LH_AOI21X2 U4316 ( .A(n6016), .B(n6083), .C(n6015), .Z(n6017) );
  HS65_LH_NAND2X4 U4317 ( .A(n8574), .B(n3407), .Z(n3344) );
  HS65_LH_NAND2X5 U4320 ( .A(n4213), .B(n7869), .Z(n8565) );
  HS65_LH_OAI12X3 U4323 ( .A(n8177), .B(n8132), .C(n2733), .Z(n8133) );
  HS65_LL_NAND2X4 U4324 ( .A(n9213), .B(n7118), .Z(n7796) );
  HS65_LH_NAND2X4 U4325 ( .A(n9112), .B(n8576), .Z(n8134) );
  HS65_LH_AOI12X2 U4326 ( .A(n5808), .B(n5868), .C(n5807), .Z(n5809) );
  HS65_LH_NAND2X5 U4327 ( .A(n3127), .B(n3407), .Z(n4971) );
  HS65_LH_OAI21X2 U4328 ( .A(n7762), .B(n7761), .C(n7760), .Z(n8124) );
  HS65_LH_NAND2X4 U4330 ( .A(n3193), .B(n7802), .Z(n8533) );
  HS65_LL_NAND2X21 U4332 ( .A(n2733), .B(n8034), .Z(
        \u_DataPath/u_fetch/pc1/N3 ) );
  HS65_LL_OAI12X3 U4333 ( .A(n5736), .B(n5799), .C(n5735), .Z(n5904) );
  HS65_LL_BFX27 U4334 ( .A(n7802), .Z(n7869) );
  HS65_LL_IVX9 U4335 ( .A(n3333), .Z(n3407) );
  HS65_LH_NOR2X5 U4336 ( .A(n7724), .B(n7720), .Z(n7721) );
  HS65_LH_NAND2X4 U4337 ( .A(n3256), .B(n7802), .Z(n8515) );
  HS65_LH_IVX7 U4338 ( .A(n2879), .Z(n3110) );
  HS65_LH_NAND2X5 U4339 ( .A(n8680), .B(n7746), .Z(n7747) );
  HS65_LH_IVX9 U4340 ( .A(n7614), .Z(n7615) );
  HS65_LH_NOR2X5 U4341 ( .A(n7834), .B(n3968), .Z(n4192) );
  HS65_LH_IVX7 U4342 ( .A(n7903), .Z(n4243) );
  HS65_LL_IVX18 U4343 ( .A(n3308), .Z(n7802) );
  HS65_LHS_XNOR2X3 U4344 ( .A(n6104), .B(n6103), .Z(
        \u_DataPath/u_execute/resAdd1_i [3]) );
  HS65_LH_IVX7 U4347 ( .A(n3111), .Z(n8577) );
  HS65_LL_NAND2X5 U4349 ( .A(n2981), .B(n3111), .Z(n3114) );
  HS65_LHS_XOR2X3 U4350 ( .A(n7788), .B(n7787), .Z(
        \u_DataPath/u_execute/link_value_i [6]) );
  HS65_LH_NOR2X5 U4351 ( .A(n5932), .B(n5964), .Z(n5934) );
  HS65_LH_NOR2X6 U4352 ( .A(n7680), .B(n7741), .Z(n7746) );
  HS65_LL_NOR2X5 U4355 ( .A(n6349), .B(n6333), .Z(n6746) );
  HS65_LH_CNIVX3 U4356 ( .A(n5798), .Z(n5802) );
  HS65_LH_IVX7 U4357 ( .A(n7676), .Z(n7678) );
  HS65_LH_CNIVX3 U4358 ( .A(n8284), .Z(\u_DataPath/branch_target_i [0]) );
  HS65_LH_NOR2X6 U4359 ( .A(n5730), .B(n5760), .Z(n5732) );
  HS65_LH_NOR3X4 U4360 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .B(n8162), 
        .C(n7703), .Z(n8098) );
  HS65_LH_NAND2X5 U4361 ( .A(n2733), .B(n8266), .Z(n8304) );
  HS65_LH_NAND2X4 U4362 ( .A(n2733), .B(n8255), .Z(n8293) );
  HS65_LH_IVX4 U4363 ( .A(n8380), .Z(n4207) );
  HS65_LH_AOI21X6 U4364 ( .A(n6051), .B(n5922), .C(n5921), .Z(n6034) );
  HS65_LH_NAND2X5 U4365 ( .A(n8316), .B(n2733), .Z(n8321) );
  HS65_LH_NAND2X5 U4368 ( .A(n2733), .B(n8243), .Z(n8362) );
  HS65_LH_NAND2X4 U4370 ( .A(n2733), .B(\u_DataPath/toPC2_i [0]), .Z(n8284) );
  HS65_LH_IVX9 U4371 ( .A(n8323), .Z(n8537) );
  HS65_LH_NAND2X5 U4372 ( .A(n2733), .B(n8176), .Z(n8422) );
  HS65_LH_NAND2X4 U4373 ( .A(n2733), .B(n8339), .Z(n8343) );
  HS65_LH_NAND2X5 U4374 ( .A(n2733), .B(n8374), .Z(n8378) );
  HS65_LH_NAND2X4 U4375 ( .A(n2733), .B(n8394), .Z(n8434) );
  HS65_LH_NAND2X5 U4376 ( .A(n2733), .B(n8364), .Z(n8367) );
  HS65_LH_NAND2X5 U4377 ( .A(n2733), .B(n8355), .Z(n8358) );
  HS65_LH_NAND2X5 U4378 ( .A(n2733), .B(n8550), .Z(n8372) );
  HS65_LH_OAI21X6 U4379 ( .A(n3404), .B(n3023), .C(n3022), .Z(n5716) );
  HS65_LH_IVX4 U4380 ( .A(n5844), .Z(n5898) );
  HS65_LH_NAND2X4 U4381 ( .A(n2733), .B(n8332), .Z(n8337) );
  HS65_LH_IVX4 U4382 ( .A(n5757), .Z(n5763) );
  HS65_LH_IVX4 U4383 ( .A(n5761), .Z(n5762) );
  HS65_LH_CNIVX3 U4385 ( .A(n5779), .Z(n5782) );
  HS65_LH_NAND2X4 U4386 ( .A(n2733), .B(n8389), .Z(n8404) );
  HS65_LH_IVX9 U4387 ( .A(n4175), .Z(n3288) );
  HS65_LH_NAND2X5 U4389 ( .A(n2733), .B(n8393), .Z(n8431) );
  HS65_LL_NOR3X2 U4391 ( .A(\u_DataPath/cw_to_ex_i [15]), .B(n8755), .C(n8263), 
        .Z(n8451) );
  HS65_LH_NOR2X2 U4393 ( .A(n8065), .B(rst), .Z(
        \u_DataPath/regfile_addr_out_towb_i [2]) );
  HS65_LH_NOR2X5 U4395 ( .A(n8042), .B(rst), .Z(\u_DataPath/idex_rt_i [3]) );
  HS65_LH_IVX4 U4397 ( .A(n5687), .Z(n5689) );
  HS65_LH_NOR2X2 U4398 ( .A(n8108), .B(rst), .Z(
        \u_DataPath/regfile_addr_out_towb_i [0]) );
  HS65_LH_NOR2X3 U4399 ( .A(n8574), .B(rst), .Z(n8579) );
  HS65_LL_NAND2X5 U4401 ( .A(\u_DataPath/jaddr_i [16]), .B(n8153), .Z(n6353)
         );
  HS65_LH_NAND2X5 U4402 ( .A(n2733), .B(n8311), .Z(n8314) );
  HS65_LH_CNIVX3 U4403 ( .A(n7725), .Z(n7789) );
  HS65_LH_NOR2X2 U4405 ( .A(n8063), .B(rst), .Z(
        \u_DataPath/regfile_addr_out_towb_i [3]) );
  HS65_LH_IVX4 U4406 ( .A(n5820), .Z(n5866) );
  HS65_LH_NAND2X2 U4407 ( .A(\u_DataPath/cw_to_ex_i [2]), .B(n7834), .Z(n4786)
         );
  HS65_LH_IVX7 U4408 ( .A(\u_DataPath/dataOut_exe_i [24]), .Z(n3140) );
  HS65_LH_IVX4 U4409 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .Z(n8130) );
  HS65_LH_IVX4 U4410 ( .A(n9077), .Z(n2943) );
  HS65_LH_NAND2X5 U4412 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [10]), 
        .Z(n8182) );
  HS65_LH_NAND2X5 U4413 ( .A(n9177), .B(n9229), .Z(n5877) );
  HS65_LH_NAND2X5 U4416 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [9]), 
        .Z(n8185) );
  HS65_LH_NAND2X5 U4417 ( .A(n9030), .B(n9223), .Z(n5838) );
  HS65_LH_NAND2X5 U4418 ( .A(n9343), .B(n9221), .Z(n5819) );
  HS65_LH_NAND2X7 U4419 ( .A(n9223), .B(n9219), .Z(n4001) );
  HS65_LH_NOR2X6 U4420 ( .A(n9341), .B(n9218), .Z(n5795) );
  HS65_LH_NAND2X2 U4421 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [2]), .Z(
        n8228) );
  HS65_LH_NAND2X2 U4422 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [0]), .Z(
        n8230) );
  HS65_LH_NAND2X5 U4424 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [8]), 
        .Z(n8186) );
  HS65_LH_IVX7 U4425 ( .A(\u_DataPath/dataOut_exe_i [18]), .Z(n3193) );
  HS65_LH_NOR2X6 U4427 ( .A(n9267), .B(n9228), .Z(n5786) );
  HS65_LH_NOR3X3 U4428 ( .A(n8755), .B(n9151), .C(\u_DataPath/cw_to_ex_i [15]), 
        .Z(n8264) );
  HS65_LH_NAND2X5 U4430 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [7]), 
        .Z(n8179) );
  HS65_LH_IVX4 U4431 ( .A(n8876), .Z(n4715) );
  HS65_LH_IVX9 U4432 ( .A(\u_DataPath/dataOut_exe_i [25]), .Z(n3132) );
  HS65_LH_NAND2X5 U4433 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [6]), 
        .Z(n8187) );
  HS65_LH_NAND2X2 U4435 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [20]), 
        .Z(n8205) );
  HS65_LH_NAND2X2 U4436 ( .A(n2733), .B(n9427), .Z(n8196) );
  HS65_LH_IVX7 U4437 ( .A(n9236), .Z(n2975) );
  HS65_LH_NAND2X2 U4438 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [6]), .Z(
        n8224) );
  HS65_LH_IVX7 U4439 ( .A(\u_DataPath/dataOut_exe_i [13]), .Z(n3252) );
  HS65_LH_IVX7 U4440 ( .A(\u_DataPath/dataOut_exe_i [4]), .Z(n8574) );
  HS65_LH_IVX9 U4441 ( .A(\u_DataPath/from_mem_data_out_i [1]), .Z(n3021) );
  HS65_LH_NAND2X2 U4442 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [19]), 
        .Z(n8206) );
  HS65_LH_NAND2X2 U4443 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [27]), 
        .Z(n8194) );
  HS65_LH_NOR2X5 U4444 ( .A(n8943), .B(n9210), .Z(n6026) );
  HS65_LH_NAND2X2 U4445 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [7]), .Z(
        n8223) );
  HS65_LH_NAND2X2 U4446 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [8]), .Z(
        n8222) );
  HS65_LH_NAND2X2 U4447 ( .A(n2733), .B(n9426), .Z(n8208) );
  HS65_LH_NAND2X2 U4448 ( .A(n2733), .B(n9425), .Z(n8193) );
  HS65_LH_NAND2X2 U4449 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [17]), 
        .Z(n8209) );
  HS65_LH_NAND2X2 U4450 ( .A(n2733), .B(n9424), .Z(n8211) );
  HS65_LH_IVX7 U4451 ( .A(\u_DataPath/dataOut_exe_i [11]), .Z(n3232) );
  HS65_LH_NAND2X2 U4452 ( .A(n2733), .B(n9423), .Z(n8221) );
  HS65_LH_NAND2X2 U4455 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [29]), 
        .Z(n8191) );
  HS65_LH_NAND2X7 U4456 ( .A(n8968), .B(n9217), .Z(n5997) );
  HS65_LH_NAND2X2 U4457 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [10]), 
        .Z(n8219) );
  HS65_LH_NAND2X7 U4458 ( .A(n9077), .B(n9218), .Z(n6063) );
  HS65_LH_NAND2X2 U4459 ( .A(n2733), .B(n9422), .Z(n8218) );
  HS65_LH_NAND2X2 U4460 ( .A(n2733), .B(n9421), .Z(n8190) );
  HS65_LH_NAND2X2 U4461 ( .A(n2733), .B(n9419), .Z(n8216) );
  HS65_LH_IVX7 U4462 ( .A(\u_DataPath/dataOut_exe_i [10]), .Z(n3242) );
  HS65_LH_NAND2X2 U4463 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [13]), 
        .Z(n8214) );
  HS65_LH_NAND2X2 U4464 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [15]), 
        .Z(n8212) );
  HS65_LH_IVX4 U4465 ( .A(n9226), .Z(n7724) );
  HS65_LH_NAND2X2 U4466 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [31]), 
        .Z(n8289) );
  HS65_LH_NAND2X2 U4467 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [14]), 
        .Z(n8213) );
  HS65_LH_NAND2X2 U4468 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [1]), .Z(
        n8229) );
  HS65_LH_IVX9 U4469 ( .A(n8724), .Z(n3345) );
  HS65_LH_NAND2X5 U4470 ( .A(n9033), .B(n9215), .Z(n6099) );
  HS65_LH_NAND2X7 U4471 ( .A(n8913), .B(n9219), .Z(n6094) );
  HS65_LH_NAND2X2 U4472 ( .A(n2733), .B(n9420), .Z(n8200) );
  HS65_LH_IVX2 U4474 ( .A(n9116), .Z(\u_DataPath/u_execute/link_value_i [2])
         );
  HS65_LH_NAND2X7 U4475 ( .A(n9030), .B(n9223), .Z(n6040) );
  HS65_LH_NAND2X2 U4476 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [3]), .Z(
        n8227) );
  HS65_LH_NAND2X2 U4477 ( .A(n2733), .B(n9429), .Z(n8202) );
  HS65_LH_NAND2X2 U4478 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [25]), 
        .Z(n8197) );
  HS65_LH_NAND2X2 U4479 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [4]), .Z(
        n8226) );
  HS65_LH_NAND2X2 U4480 ( .A(n2733), .B(n9428), .Z(n8204) );
  HS65_LH_IVX4 U4481 ( .A(n9230), .Z(n7793) );
  HS65_LH_NAND2X2 U4483 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [5]), .Z(
        n8225) );
  HS65_LH_NAND2X2 U4484 ( .A(n2733), .B(\u_DataPath/pc4_to_idexreg_i [24]), 
        .Z(n8198) );
  HS65_LH_IVX7 U4487 ( .A(\u_DataPath/dataOut_exe_i [5]), .Z(n3336) );
  HS65_LL_IVX7 U4489 ( .A(\u_DataPath/jaddr_i [16]), .Z(n8152) );
  HS65_LH_IVX2 U4490 ( .A(Data_out_fromRAM[30]), .Z(n8402) );
  HS65_LH_IVX2 U4491 ( .A(Data_out_fromRAM[29]), .Z(n8447) );
  HS65_LH_IVX2 U4493 ( .A(Data_out_fromRAM[24]), .Z(n8370) );
  HS65_LH_IVX2 U4494 ( .A(Data_out_fromRAM[27]), .Z(n8376) );
  HS65_LH_IVX2 U4495 ( .A(Data_out_fromRAM[26]), .Z(n8319) );
  HS65_LH_IVX2 U4496 ( .A(Data_out_fromRAM[25]), .Z(n8335) );
  HS65_LH_OAI12X6 U4497 ( .A(n5715), .B(n5714), .C(n5713), .Z(n7860) );
  HS65_LL_NAND2X4 U4498 ( .A(n7907), .B(n5694), .Z(n7855) );
  HS65_LL_NAND2X2 U4499 ( .A(n7858), .B(n9063), .Z(
        \u_DataPath/dataOut_exe_i [19]) );
  HS65_LL_OAI12X3 U4501 ( .A(n9189), .B(n9001), .C(n8395), .Z(
        \u_DataPath/dataOut_exe_i [30]) );
  HS65_LL_OAI12X3 U4502 ( .A(n9189), .B(n8895), .C(n8398), .Z(
        \u_DataPath/dataOut_exe_i [14]) );
  HS65_LL_NAND2X2 U4503 ( .A(n7845), .B(n9060), .Z(
        \u_DataPath/dataOut_exe_i [21]) );
  HS65_LL_OAI12X3 U4505 ( .A(n9189), .B(n8889), .C(n8405), .Z(
        \u_DataPath/dataOut_exe_i [17]) );
  HS65_LL_AOI21X2 U4508 ( .A(n5643), .B(n5642), .C(n5641), .Z(n5674) );
  HS65_LH_NAND2X7 U4509 ( .A(n7843), .B(n9062), .Z(
        \u_DataPath/dataOut_exe_i [18]) );
  HS65_LL_OAI12X3 U4510 ( .A(n9189), .B(n9059), .C(n8409), .Z(
        \u_DataPath/dataOut_exe_i [20]) );
  HS65_LL_NOR2AX3 U4511 ( .A(n4912), .B(n4911), .Z(n8474) );
  HS65_LL_NAND2X2 U4512 ( .A(n4910), .B(n4909), .Z(n4911) );
  HS65_LL_NAND2X2 U4513 ( .A(n3695), .B(n3694), .Z(n3696) );
  HS65_LH_AOI21X6 U4514 ( .A(n5643), .B(n4280), .C(n4279), .Z(n4281) );
  HS65_LH_NAND2X7 U4515 ( .A(n5643), .B(n3624), .Z(n3625) );
  HS65_LH_NAND2X7 U4518 ( .A(n5643), .B(n3742), .Z(n3743) );
  HS65_LL_NAND3X3 U4519 ( .A(n3998), .B(n3997), .C(n3996), .Z(n3999) );
  HS65_LH_NAND2X7 U4520 ( .A(n5643), .B(n3693), .Z(n3694) );
  HS65_LHS_XNOR2X6 U4521 ( .A(n4429), .B(n4428), .Z(n4450) );
  HS65_LL_OAI21X2 U4522 ( .A(n5633), .B(n4240), .C(n4239), .Z(n4241) );
  HS65_LH_AOI21X6 U4523 ( .A(n5285), .B(n4569), .C(n4568), .Z(n8464) );
  HS65_LH_OAI12X3 U4524 ( .A(n4377), .B(n2859), .C(n4376), .Z(n4378) );
  HS65_LL_OAI21X2 U4525 ( .A(n2859), .B(n3739), .C(n3738), .Z(n3740) );
  HS65_LH_OAI12X3 U4527 ( .A(n3706), .B(n5633), .C(n3705), .Z(n3707) );
  HS65_LHS_XOR2X3 U4529 ( .A(n4847), .B(n2859), .Z(n4861) );
  HS65_LH_NOR2AX3 U4530 ( .A(n5672), .B(n5251), .Z(n5252) );
  HS65_LL_OAI21X2 U4531 ( .A(n2859), .B(n4224), .C(n4223), .Z(n4225) );
  HS65_LL_OAI21X2 U4532 ( .A(n3621), .B(n2859), .C(n3620), .Z(n3622) );
  HS65_LH_AOI21X6 U4533 ( .A(n5285), .B(n4605), .C(n4604), .Z(n8463) );
  HS65_LH_AOI12X2 U4534 ( .A(n3634), .B(n5195), .C(n3633), .Z(n3635) );
  HS65_LH_OAI21X3 U4535 ( .A(n4993), .B(n4992), .C(n4991), .Z(n4994) );
  HS65_LH_IVX4 U4536 ( .A(n4473), .Z(n4446) );
  HS65_LL_AOI21X2 U4537 ( .A(n5492), .B(n4781), .C(n5122), .Z(n5159) );
  HS65_LH_IVX4 U4538 ( .A(n5559), .Z(n5539) );
  HS65_LH_IVX4 U4539 ( .A(n5210), .Z(n5213) );
  HS65_LH_NAND2X5 U4541 ( .A(n3688), .B(n5210), .Z(n3690) );
  HS65_LH_NAND3X3 U4543 ( .A(n5515), .B(n4050), .C(n5526), .Z(n5110) );
  HS65_LH_OAI21X3 U4546 ( .A(n4751), .B(n5656), .C(n3771), .Z(n3787) );
  HS65_LL_OAI12X3 U4550 ( .A(n4085), .B(n3481), .C(n3479), .Z(n3617) );
  HS65_LH_NAND2X4 U4551 ( .A(n4222), .B(n5210), .Z(n4224) );
  HS65_LH_NAND2X4 U4552 ( .A(n5429), .B(n5458), .Z(n5461) );
  HS65_LH_NAND2X4 U4553 ( .A(n5029), .B(n5028), .Z(n5076) );
  HS65_LH_NAND2X4 U4555 ( .A(n4528), .B(n4164), .Z(n3767) );
  HS65_LL_IVX4 U4558 ( .A(n4928), .Z(n4085) );
  HS65_LH_NAND2X4 U4560 ( .A(n3737), .B(n2867), .Z(n3739) );
  HS65_LH_NAND2X4 U4562 ( .A(n3704), .B(n5631), .Z(n3706) );
  HS65_LH_NAND2X5 U4563 ( .A(n4916), .B(n3897), .Z(n3899) );
  HS65_LH_NAND2X4 U4564 ( .A(n5131), .B(n4578), .Z(n3914) );
  HS65_LH_NAND2AX7 U4565 ( .A(n4689), .B(n4688), .Z(n4693) );
  HS65_LH_OAI12X3 U4566 ( .A(n5147), .B(n5146), .C(n5145), .Z(n5148) );
  HS65_LH_NAND2X7 U4567 ( .A(n5488), .B(n5487), .Z(n5489) );
  HS65_LH_NAND3X5 U4568 ( .A(n4757), .B(n4945), .C(n4756), .Z(n4758) );
  HS65_LH_IVX9 U4569 ( .A(n4522), .Z(n5666) );
  HS65_LH_NAND2X4 U4570 ( .A(n4396), .B(n4395), .Z(n4397) );
  HS65_LH_NOR2X6 U4571 ( .A(n4913), .B(n3282), .Z(n3897) );
  HS65_LH_OAI12X3 U4572 ( .A(n5456), .B(n5455), .C(n5454), .Z(n5457) );
  HS65_LH_NOR2X5 U4574 ( .A(n5456), .B(n5428), .Z(n5458) );
  HS65_LH_NOR2X3 U4575 ( .A(n4955), .B(n5146), .Z(n4956) );
  HS65_LH_OAI211X4 U4577 ( .A(n5656), .B(n4613), .C(n4612), .D(n4611), .Z(
        n4620) );
  HS65_LH_OAI21X3 U4579 ( .A(n5412), .B(n5411), .C(n5410), .Z(n5413) );
  HS65_LH_NOR2X3 U4580 ( .A(n5646), .B(n4119), .Z(n4123) );
  HS65_LH_NOR2X5 U4581 ( .A(n4220), .B(n4317), .Z(n4222) );
  HS65_LH_NAND2X5 U4582 ( .A(n5661), .B(n5174), .Z(n5175) );
  HS65_LH_AOI12X2 U4583 ( .A(n4476), .B(n4632), .C(n4109), .Z(n4110) );
  HS65_LH_IVX7 U4584 ( .A(n4391), .Z(n3522) );
  HS65_LH_IVX7 U4586 ( .A(n4291), .Z(n4292) );
  HS65_LH_NAND3X3 U4587 ( .A(n5237), .B(n5236), .C(n5235), .Z(n5238) );
  HS65_LH_NAND2X5 U4588 ( .A(n3792), .B(n3791), .Z(n3793) );
  HS65_LH_OAI21X3 U4589 ( .A(n5646), .B(n4522), .C(n4267), .Z(n4275) );
  HS65_LH_IVX9 U4590 ( .A(n3913), .Z(n4578) );
  HS65_LH_NOR3X4 U4591 ( .A(n4710), .B(n4730), .C(n4709), .Z(n4733) );
  HS65_LH_NAND2X5 U4592 ( .A(n5643), .B(n4599), .Z(n4600) );
  HS65_LH_IVX7 U4593 ( .A(n4332), .Z(n3388) );
  HS65_LH_AOI22X4 U4594 ( .A(n5131), .B(n4157), .C(n4887), .D(n4950), .Z(n4171) );
  HS65_LH_NAND2X4 U4595 ( .A(n5661), .B(n5203), .Z(n3461) );
  HS65_LH_NAND2X4 U4597 ( .A(n5618), .B(n5243), .Z(n3712) );
  HS65_LH_IVX4 U4598 ( .A(n4185), .Z(n3723) );
  HS65_LH_NOR2X6 U4599 ( .A(n5510), .B(n5583), .Z(n5536) );
  HS65_LH_IVX9 U4604 ( .A(n4176), .Z(n5240) );
  HS65_LH_IVX7 U4605 ( .A(n5505), .Z(n5562) );
  HS65_LH_IVX9 U4608 ( .A(n4393), .Z(n4889) );
  HS65_LH_NOR2X5 U4609 ( .A(n4320), .B(n4317), .Z(n4322) );
  HS65_LH_NOR2X3 U4610 ( .A(n4333), .B(n4330), .Z(n4335) );
  HS65_LH_AOI22X3 U4612 ( .A(n4508), .B(n4344), .C(n4516), .D(n4120), .Z(n3557) );
  HS65_LH_NAND2X7 U4613 ( .A(n4015), .B(n4017), .Z(n3952) );
  HS65_LH_IVX7 U4615 ( .A(n4290), .Z(n4293) );
  HS65_LH_NOR2X5 U4617 ( .A(n3800), .B(n3685), .Z(n3688) );
  HS65_LH_IVX9 U4618 ( .A(n3905), .Z(n4007) );
  HS65_LH_NOR2X5 U4621 ( .A(n3747), .B(n3631), .Z(n3634) );
  HS65_LH_NAND3X3 U4622 ( .A(n4672), .B(n5517), .C(n5296), .Z(n5333) );
  HS65_LL_AOI21X2 U4623 ( .A(n5208), .B(n5211), .C(n3619), .Z(n3620) );
  HS65_LH_NAND2X5 U4624 ( .A(n5453), .B(n5424), .Z(n5456) );
  HS65_LH_NOR3X3 U4626 ( .A(n5522), .B(n5542), .C(n5099), .Z(n5100) );
  HS65_LH_NAND2X5 U4627 ( .A(n4774), .B(n4773), .Z(n4775) );
  HS65_LH_IVX9 U4628 ( .A(n4317), .Z(n3505) );
  HS65_LH_OAI21X3 U4630 ( .A(n3863), .B(n3862), .C(n5229), .Z(n3864) );
  HS65_LH_OAI211X3 U4631 ( .A(n5360), .B(n5359), .C(n5358), .D(n5478), .Z(
        n5369) );
  HS65_LH_NAND2X7 U4632 ( .A(n3574), .B(n3573), .Z(n3580) );
  HS65_LH_CNIVX3 U4635 ( .A(n3375), .Z(n3210) );
  HS65_LH_NAND2X4 U4636 ( .A(n5446), .B(n5427), .Z(n5428) );
  HS65_LH_NAND2X5 U4639 ( .A(n3684), .B(n3683), .Z(n3692) );
  HS65_LH_IVX7 U4640 ( .A(n4038), .Z(n4039) );
  HS65_LH_NAND3X5 U4641 ( .A(n4591), .B(n4590), .C(n4589), .Z(n4617) );
  HS65_LH_IVX9 U4642 ( .A(n4426), .Z(n5607) );
  HS65_LH_IVX9 U4644 ( .A(n4835), .Z(n4468) );
  HS65_LH_AOI22X3 U4645 ( .A(n9349), .B(n5321), .C(n5131), .D(n4584), .Z(n4585) );
  HS65_LH_IVX4 U4646 ( .A(n4894), .Z(n3598) );
  HS65_LH_AOI12X2 U4647 ( .A(n3586), .B(n3585), .C(n4581), .Z(n3588) );
  HS65_LH_NAND3X3 U4648 ( .A(n5469), .B(n5468), .C(n5467), .Z(n5470) );
  HS65_LH_NOR2X3 U4649 ( .A(n4643), .B(n4639), .Z(n4646) );
  HS65_LH_NAND2X7 U4650 ( .A(n3650), .B(n3649), .Z(n3651) );
  HS65_LH_IVX4 U4651 ( .A(n4496), .Z(n4499) );
  HS65_LH_OA12X9 U4652 ( .A(n5656), .B(n4945), .C(n4944), .Z(n2898) );
  HS65_LH_AOI12X2 U4654 ( .A(n5139), .B(n5229), .C(n5138), .Z(n5140) );
  HS65_LH_NOR2X3 U4655 ( .A(n4134), .B(n4939), .Z(n4610) );
  HS65_LH_NOR2X5 U4656 ( .A(n5627), .B(n3701), .Z(n3704) );
  HS65_LH_IVX7 U4657 ( .A(n5499), .Z(n5563) );
  HS65_LH_NAND2X4 U4658 ( .A(n5547), .B(n5091), .Z(n5474) );
  HS65_LH_NOR3X4 U4660 ( .A(n4772), .B(n4771), .C(n4770), .Z(n4773) );
  HS65_LH_NOR2X3 U4661 ( .A(n4328), .B(n4333), .Z(n5424) );
  HS65_LH_NAND2X7 U4662 ( .A(n3615), .B(n3614), .Z(n3623) );
  HS65_LH_NAND2X5 U4663 ( .A(n3750), .B(n3383), .Z(n3387) );
  HS65_LH_NOR2X6 U4664 ( .A(n3640), .B(n3639), .Z(n3643) );
  HS65_LH_NOR2X5 U4666 ( .A(n5389), .B(n4667), .Z(n4668) );
  HS65_LH_NAND2X7 U4667 ( .A(n4154), .B(n3867), .Z(n3863) );
  HS65_LH_IVX4 U4668 ( .A(n5514), .Z(n5520) );
  HS65_LH_NAND2X7 U4669 ( .A(n4542), .B(n4462), .Z(n3862) );
  HS65_LH_IVX7 U4670 ( .A(n5083), .Z(n5304) );
  HS65_LH_NAND2X7 U4671 ( .A(n5344), .B(n5564), .Z(n4720) );
  HS65_LH_OAI12X3 U4672 ( .A(n5183), .B(n5182), .C(n5181), .Z(n5184) );
  HS65_LH_IVX4 U4673 ( .A(n4580), .Z(n4552) );
  HS65_LH_IVX4 U4675 ( .A(n5545), .Z(n5557) );
  HS65_LH_NAND2X5 U4676 ( .A(n3529), .B(n3444), .Z(n4488) );
  HS65_LH_NOR2X6 U4677 ( .A(n5363), .B(n5471), .Z(n5507) );
  HS65_LH_NAND2X4 U4679 ( .A(n5300), .B(n5516), .Z(n5479) );
  HS65_LH_NAND2X4 U4680 ( .A(n5357), .B(n5356), .Z(n5478) );
  HS65_LH_NOR2X6 U4681 ( .A(n4984), .B(n4582), .Z(n3982) );
  HS65_LH_IVX4 U4682 ( .A(n4462), .Z(n4464) );
  HS65_LH_IVX4 U4683 ( .A(n4059), .Z(n3535) );
  HS65_LH_OAI12X3 U4684 ( .A(n2848), .B(n4795), .C(n3524), .Z(n3528) );
  HS65_LH_IVX7 U4686 ( .A(n4027), .Z(n4031) );
  HS65_LH_NAND2X5 U4687 ( .A(n3749), .B(n3748), .Z(n3755) );
  HS65_LH_IVX7 U4688 ( .A(n3867), .Z(n3868) );
  HS65_LH_IVX7 U4689 ( .A(n4289), .Z(n4218) );
  HS65_LH_IVX4 U4690 ( .A(n3956), .Z(n3957) );
  HS65_LH_NAND2X5 U4692 ( .A(n5531), .B(n5293), .Z(n3517) );
  HS65_LH_IVX9 U4693 ( .A(n5571), .Z(n4727) );
  HS65_LH_NAND2X7 U4694 ( .A(n3544), .B(n3543), .Z(n3546) );
  HS65_LH_NAND2X4 U4695 ( .A(n5534), .B(n5356), .Z(n5360) );
  HS65_LH_IVX4 U4696 ( .A(n5500), .Z(n5501) );
  HS65_LH_NAND2X4 U4698 ( .A(n5437), .B(n5420), .Z(n5441) );
  HS65_LH_NAND2X5 U4699 ( .A(n4060), .B(n4059), .Z(n4064) );
  HS65_LH_OAI21X3 U4700 ( .A(n3756), .B(n2854), .C(n3758), .Z(n4255) );
  HS65_LH_NAND3X5 U4702 ( .A(n5232), .B(n4808), .C(n4739), .Z(n4746) );
  HS65_LH_NAND2X5 U4703 ( .A(n4062), .B(n4061), .Z(n4063) );
  HS65_LH_IVX4 U4704 ( .A(n3682), .Z(n3683) );
  HS65_LH_NOR2X6 U4706 ( .A(n4811), .B(n4582), .Z(n3400) );
  HS65_LH_IVX9 U4709 ( .A(n5450), .Z(n4231) );
  HS65_LH_IVX9 U4710 ( .A(n5183), .Z(n5139) );
  HS65_LH_IVX7 U4711 ( .A(n4022), .Z(n4024) );
  HS65_LH_IVX4 U4714 ( .A(n5502), .Z(n5012) );
  HS65_LH_NAND2X4 U4716 ( .A(\sub_x_53/A[29] ), .B(n4587), .Z(n3441) );
  HS65_LH_NAND2X7 U4717 ( .A(n5387), .B(n5324), .Z(n5464) );
  HS65_LH_IVX4 U4718 ( .A(n4340), .Z(n4066) );
  HS65_LH_NAND2X7 U4719 ( .A(n2854), .B(n5567), .Z(n5344) );
  HS65_LH_IVX9 U4720 ( .A(n4374), .Z(n4424) );
  HS65_LH_IVX9 U4721 ( .A(n4627), .Z(n4629) );
  HS65_LH_NOR2X6 U4722 ( .A(\sub_x_53/A[29] ), .B(n5447), .Z(n4328) );
  HS65_LH_NAND2X5 U4724 ( .A(n5509), .B(n5508), .Z(n5583) );
  HS65_LH_NOR2AX3 U4725 ( .A(n5136), .B(\sub_x_53/A[0] ), .Z(n5035) );
  HS65_LH_NAND2X4 U4726 ( .A(n4628), .B(n4158), .Z(n4160) );
  HS65_LH_NAND2X7 U4727 ( .A(\lte_x_59/B[1] ), .B(n4587), .Z(n5128) );
  HS65_LH_NAND2X5 U4728 ( .A(n4819), .B(n4818), .Z(n4820) );
  HS65_LH_NAND2X4 U4729 ( .A(\sub_x_53/A[30] ), .B(n2873), .Z(n5450) );
  HS65_LH_NAND2X5 U4730 ( .A(n5098), .B(n5552), .Z(n5556) );
  HS65_LH_IVX7 U4731 ( .A(n4425), .Z(n4375) );
  HS65_LH_NAND2X5 U4732 ( .A(n5097), .B(n5096), .Z(n5545) );
  HS65_LH_NAND2X5 U4733 ( .A(\lte_x_59/B[24] ), .B(n4544), .Z(n3964) );
  HS65_LH_NOR2X3 U4734 ( .A(n3698), .B(n5627), .Z(n5437) );
  HS65_LH_NOR2X6 U4735 ( .A(n4675), .B(n4674), .Z(n5514) );
  HS65_LH_CNIVX3 U4736 ( .A(n4407), .Z(n4408) );
  HS65_LH_IVX7 U4737 ( .A(n4846), .Z(n3561) );
  HS65_LH_NAND2X7 U4738 ( .A(\sub_x_53/A[27] ), .B(n2845), .Z(n3758) );
  HS65_LL_NOR2X2 U4739 ( .A(n5254), .B(n4250), .Z(n3497) );
  HS65_LHS_XOR2X3 U4740 ( .A(n5747), .B(n5746), .Z(\u_DataPath/toPC2_i [28])
         );
  HS65_LH_IVX9 U4741 ( .A(n5530), .Z(n5295) );
  HS65_LH_NOR2X6 U4743 ( .A(n4144), .B(n4100), .Z(n4638) );
  HS65_LH_IVX9 U4745 ( .A(n3641), .Z(n4794) );
  HS65_LL_NAND2X4 U4746 ( .A(\sub_x_53/A[25] ), .B(n3593), .Z(n3615) );
  HS65_LH_IVX9 U4747 ( .A(\sub_x_53/A[0] ), .Z(n4660) );
  HS65_LH_NOR2X6 U4748 ( .A(\sub_x_53/A[25] ), .B(n3593), .Z(n3613) );
  HS65_LH_IVX9 U4749 ( .A(n4144), .Z(n4099) );
  HS65_LH_IVX9 U4750 ( .A(n3558), .Z(n3472) );
  HS65_LH_IVX4 U4751 ( .A(n3893), .Z(n4678) );
  HS65_LH_NAND2X5 U4752 ( .A(\sub_x_53/A[27] ), .B(n4588), .Z(n3650) );
  HS65_LH_NOR2X6 U4753 ( .A(\sub_x_53/A[0] ), .B(n5123), .Z(n4821) );
  HS65_LH_IVX9 U4754 ( .A(n3616), .Z(n5208) );
  HS65_LL_IVX4 U4756 ( .A(n4516), .Z(n4842) );
  HS65_LL_NAND2X4 U4757 ( .A(n3236), .B(n3238), .Z(n3239) );
  HS65_LH_IVX9 U4759 ( .A(\lte_x_59/B[21] ), .Z(n4701) );
  HS65_LH_NOR2X6 U4760 ( .A(n2858), .B(n5398), .Z(n4011) );
  HS65_LH_NAND2X7 U4761 ( .A(\lte_x_59/B[9] ), .B(n2871), .Z(n4904) );
  HS65_LH_NOR2X6 U4763 ( .A(\lte_x_59/B[22] ), .B(n2869), .Z(n5627) );
  HS65_LH_NAND3X3 U4765 ( .A(n2851), .B(n5136), .C(n4805), .Z(n4340) );
  HS65_LH_NOR2X6 U4766 ( .A(\sub_x_53/A[20] ), .B(n4699), .Z(n4374) );
  HS65_LH_NOR2X5 U4767 ( .A(\lte_x_59/B[15] ), .B(n4677), .Z(n5406) );
  HS65_LH_IVX4 U4769 ( .A(n5361), .Z(n5508) );
  HS65_LH_IVX4 U4770 ( .A(\lte_x_59/B[14] ), .Z(n4676) );
  HS65_LL_OAI21X2 U4772 ( .A(n4105), .B(n4477), .C(n4107), .Z(n4627) );
  HS65_LH_IVX4 U4773 ( .A(n4817), .Z(n4818) );
  HS65_LH_IVX9 U4774 ( .A(\lte_x_59/B[18] ), .Z(n4986) );
  HS65_LH_NAND2X7 U4775 ( .A(n4477), .B(n4476), .Z(n4478) );
  HS65_LH_NAND2X7 U4776 ( .A(\sub_x_53/A[17] ), .B(n5001), .Z(n3559) );
  HS65_LH_NAND2X7 U4777 ( .A(n4481), .B(n4480), .Z(n4482) );
  HS65_LH_NAND2X4 U4778 ( .A(n5234), .B(n4553), .Z(n4554) );
  HS65_LH_OAI22X3 U4779 ( .A(n8906), .B(n9186), .C(n9140), .D(n8759), .Z(
        \u_DataPath/data_read_ex_1_i [10]) );
  HS65_LH_OAI22X3 U4781 ( .A(n7306), .B(n8168), .C(n7914), .D(n8167), .Z(
        \u_DataPath/data_read_ex_1_i [1]) );
  HS65_LH_OAI22X3 U4782 ( .A(n7306), .B(n8275), .C(n7914), .D(n8274), .Z(
        \u_DataPath/data_read_ex_1_i [8]) );
  HS65_LH_OAI22X3 U4783 ( .A(n7306), .B(n8321), .C(n7914), .D(n8320), .Z(
        \u_DataPath/data_read_ex_1_i [26]) );
  HS65_LH_OAI22X3 U4784 ( .A(n7306), .B(n8434), .C(n7914), .D(n8174), .Z(
        \u_DataPath/data_read_ex_1_i [3]) );
  HS65_LH_OAI22X3 U4785 ( .A(n7306), .B(n8314), .C(n7914), .D(n8313), .Z(
        \u_DataPath/data_read_ex_1_i [6]) );
  HS65_LH_OAI22X3 U4787 ( .A(n7306), .B(n8293), .C(n7914), .D(n8292), .Z(
        \u_DataPath/data_read_ex_1_i [12]) );
  HS65_LH_OAI22X3 U4788 ( .A(n7306), .B(n8304), .C(n7914), .D(n8303), .Z(
        \u_DataPath/data_read_ex_1_i [7]) );
  HS65_LH_OAI22X3 U4789 ( .A(n7306), .B(n8326), .C(n7914), .D(n8325), .Z(
        \u_DataPath/data_read_ex_1_i [19]) );
  HS65_LH_IVX18 U4790 ( .A(n4683), .Z(n5398) );
  HS65_LH_IVX9 U4791 ( .A(n4823), .Z(n3486) );
  HS65_LH_NAND2X7 U4793 ( .A(n8258), .B(n3237), .Z(n3238) );
  HS65_LH_IVX4 U4794 ( .A(n4763), .Z(n4592) );
  HS65_LH_NOR2X5 U4795 ( .A(n5656), .B(n4762), .Z(n3879) );
  HS65_LL_NOR2X6 U4796 ( .A(n3159), .B(n3158), .Z(\sub_x_53/A[23] ) );
  HS65_LH_IVX7 U4797 ( .A(n4637), .Z(n3330) );
  HS65_LH_IVX9 U4798 ( .A(n4100), .Z(n4480) );
  HS65_LH_IVX9 U4800 ( .A(n4481), .Z(n4102) );
  HS65_LL_NOR2X3 U4802 ( .A(n3108), .B(n3107), .Z(n3547) );
  HS65_LH_OAI22X6 U4803 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [23]), .C(
        n8243), .D(n3409), .Z(n3158) );
  HS65_LL_OAI12X6 U4804 ( .A(n3173), .B(n2905), .C(n3172), .Z(n5654) );
  HS65_LL_IVX7 U4805 ( .A(n3401), .Z(n3399) );
  HS65_LH_NAND2X5 U4806 ( .A(\sub_x_53/A[2] ), .B(n5088), .Z(n4595) );
  HS65_LH_IVX4 U4807 ( .A(n8563), .Z(\u_DataPath/mem_writedata_out_i [28]) );
  HS65_LH_IVX9 U4809 ( .A(n5231), .Z(n3372) );
  HS65_LL_OAI12X3 U4810 ( .A(n7854), .B(n3409), .C(n3198), .Z(n3199) );
  HS65_LH_IVX9 U4811 ( .A(n5422), .Z(n5447) );
  HS65_LL_AOI12X4 U4812 ( .A(n6113), .B(n6115), .C(n5942), .Z(n5955) );
  HS65_LL_IVX27 U4813 ( .A(n3270), .Z(n3409) );
  HS65_LL_NAND2X2 U4815 ( .A(n3251), .B(n8517), .Z(n3255) );
  HS65_LH_NAND3X3 U4816 ( .A(n8562), .B(n8566), .C(n8561), .Z(n8563) );
  HS65_LL_NOR2X6 U4818 ( .A(n7799), .B(n7798), .Z(n7122) );
  HS65_LH_AOI22X3 U4819 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ), .D(
        n6363), .Z(n6287) );
  HS65_LH_AOI22X3 U4821 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ), .D(
        n6624), .Z(n7150) );
  HS65_LH_AO22X9 U4822 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ), .D(
        n7282), .Z(n6526) );
  HS65_LH_AOI22X3 U4823 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ), .D(
        n6624), .Z(n6292) );
  HS65_LH_AO22X9 U4824 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ), .D(
        n7282), .Z(n6446) );
  HS65_LH_AOI22X3 U4825 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ), .Z(n6800)
         );
  HS65_LH_AOI22X3 U4826 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ), .D(
        n7171), .Z(n6402) );
  HS65_LH_AOI22X3 U4827 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ), .D(
        n6624), .Z(n6272) );
  HS65_LH_AOI22X3 U4828 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ), .D(n7516), 
        .Z(n7521) );
  HS65_LH_AOI22X3 U4829 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ), .Z(n6779)
         );
  HS65_LH_AO22X9 U4830 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ), .Z(n7512)
         );
  HS65_LH_AOI22X3 U4834 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ), .D(n6384), .Z(n6643) );
  HS65_LH_AOI22X3 U4835 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ), .D(
        n7285), .Z(n6294) );
  HS65_LH_AOI22X3 U4836 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ), .D(
        n7285), .Z(n7288) );
  HS65_LH_AOI22X3 U4838 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][22] ), .D(
        n6363), .Z(n6267) );
  HS65_LH_AOI22X3 U4839 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][30] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ), .D(
        n6624), .Z(n6137) );
  HS65_LH_AO22X9 U4840 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ), .D(
        n7282), .Z(n6918) );
  HS65_LH_AO22X9 U4841 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ), .Z(n7533)
         );
  HS65_LH_AOI22X3 U4844 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ), .D(
        n7285), .Z(n6142) );
  HS65_LH_AO22X9 U4845 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ), .Z(n7487)
         );
  HS65_LH_AOI22X3 U4847 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ), .D(
        n7171), .Z(n6141) );
  HS65_LH_AOI22X3 U4849 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ), .Z(n6780)
         );
  HS65_LH_AOI22X3 U4850 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ), .D(
        n6384), .Z(n6155) );
  HS65_LH_AOI22X3 U4851 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ), .D(
        n7171), .Z(n6293) );
  HS65_LH_AOI22X3 U4852 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ), .D(n7516), 
        .Z(n6834) );
  HS65_LH_AO22X9 U4853 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ), .B(n7580), 
        .C(n7579), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ), .Z(n7387) );
  HS65_LH_AO22X9 U4854 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ), .D(
        n7282), .Z(n6381) );
  HS65_LH_AO22X9 U4856 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ), .Z(n7447)
         );
  HS65_LH_AO22X9 U4857 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ), .B(n7429), 
        .C(n6952), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ), .Z(n7388) );
  HS65_LH_AOI22X3 U4858 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ), .D(n6740), 
        .Z(n7389) );
  HS65_LH_AO22X9 U4859 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ), .Z(n7492)
         );
  HS65_LH_AOI22X3 U4861 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ), .D(
        n2888), .Z(n6227) );
  HS65_LH_AOI22X3 U4862 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][16] ), .D(
        n6624), .Z(n6170) );
  HS65_LH_AO22X9 U4865 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ), .Z(n7608)
         );
  HS65_LH_AO22X9 U4866 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ), .D(
        n6637), .Z(n6235) );
  HS65_LH_AO22X9 U4867 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ), .B(n7522), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ), .Z(n7398)
         );
  HS65_LH_AO22X9 U4869 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ), .D(
        n7292), .Z(n6239) );
  HS65_LH_AO22X9 U4871 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ), .Z(n7507)
         );
  HS65_LH_AOI22X3 U4873 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ), .D(
        n6670), .Z(n7227) );
  HS65_LH_AO22X9 U4875 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ), .Z(n7573)
         );
  HS65_LH_AO22X9 U4876 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ), .Z(n7446)
         );
  HS65_LH_AOI22X3 U4879 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ), .D(
        n6624), .Z(n6232) );
  HS65_LH_AOI22X3 U4881 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ), .Z(n7335)
         );
  HS65_LH_AO22X9 U4882 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ), .B(n7429), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ), .Z(n7493)
         );
  HS65_LH_AOI22X3 U4883 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ), .Z(n6799)
         );
  HS65_LH_AO22X9 U4884 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ), .B(n7580), 
        .C(n7579), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ), .Z(n7430) );
  HS65_LH_AOI22X3 U4885 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ), .D(n7516), 
        .Z(n6706) );
  HS65_LH_AO22X9 U4887 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ), .Z(n7553)
         );
  HS65_LH_AOI22X3 U4890 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ), .Z(n7336)
         );
  HS65_LH_AOI22X3 U4891 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ), .D(n6740), 
        .Z(n7494) );
  HS65_LH_AOI22X3 U4892 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][21] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ), .D(
        n6625), .Z(n6191) );
  HS65_LH_AOI22X3 U4893 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][5] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ), .D(n6942), .Z(n6943) );
  HS65_LH_AO22X9 U4899 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ), .Z(n7506)
         );
  HS65_LH_AOI22X3 U4900 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ), .D(n2889), .Z(n7437) );
  HS65_LH_AOI22X3 U4901 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][27] ), .D(
        n6624), .Z(n6212) );
  HS65_LH_AOI22X3 U4903 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ), .D(n7516), 
        .Z(n7499) );
  HS65_LH_AOI22X3 U4904 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ), .D(
        n7171), .Z(n6273) );
  HS65_LH_AOI22X3 U4907 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ), .D(
        n6624), .Z(n6252) );
  HS65_LH_AO22X9 U4908 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ), .Z(n7558)
         );
  HS65_LH_AOI22X3 U4910 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][11] ), .D(
        n6363), .Z(n6247) );
  HS65_LH_AOI22X3 U4911 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ), .D(
        n7171), .Z(n7172) );
  HS65_LH_AOI22X3 U4912 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ), .D(
        n2888), .Z(n6622) );
  HS65_LH_AOI22X3 U4913 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ), .D(
        n7285), .Z(n7173) );
  HS65_LH_AOI22X3 U4914 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ), .D(n7516), 
        .Z(n6679) );
  HS65_LH_AO22X9 U4916 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][11] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ), .D(
        n7292), .Z(n6259) );
  HS65_LH_AO22X9 U4918 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ), .D(
        n6637), .Z(n6255) );
  HS65_LH_AO22X9 U4919 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ), .D(
        n7282), .Z(n6425) );
  HS65_LH_AOI22X3 U4920 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ), .D(
        n6363), .Z(n7163) );
  HS65_LH_AOI22X3 U4922 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ), .D(
        n7171), .Z(n6313) );
  HS65_LH_AOI22X3 U4924 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ), .Z(n7256)
         );
  HS65_LH_AOI22X3 U4926 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ), .D(n7516), 
        .Z(n6794) );
  HS65_LH_AO22X9 U4929 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ), .Z(n7367)
         );
  HS65_LH_AOI22X3 U4930 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ), .Z(n7257)
         );
  HS65_LH_AO22X9 U4931 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ), .D(
        n6637), .Z(n6315) );
  HS65_LH_AOI22X3 U4932 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ), .D(n7516), 
        .Z(n7374) );
  HS65_LH_AOI22X3 U4935 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ), .Z(n7196)
         );
  HS65_LH_AO22X9 U4937 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ), .Z(n7467)
         );
  HS65_LH_AOI22X3 U4939 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ), .Z(n7197)
         );
  HS65_LH_AO22X9 U4940 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ), .D(
        n6637), .Z(n7133) );
  HS65_LH_AOI22X3 U4941 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ), .D(
        n6624), .Z(n6312) );
  HS65_LH_AOI22X3 U4943 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ), .D(
        n7285), .Z(n6274) );
  HS65_LH_AOI22X3 U4946 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ), .D(n7516), 
        .Z(n6814) );
  HS65_LH_AO22X9 U4947 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ), .D(
        n7282), .Z(n6405) );
  HS65_LH_AOI22X3 U4950 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ), .Z(n6796)
         );
  HS65_LH_AOI22X3 U4952 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][17] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ), .D(
        n6942), .Z(n6899) );
  HS65_LH_AO22X9 U4953 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ), .D(
        n7282), .Z(n6858) );
  HS65_LH_AOI22X3 U4954 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ), .D(
        n7264), .Z(n7271) );
  HS65_LH_AOI22X3 U4955 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ), .D(
        n6363), .Z(n7270) );
  HS65_LH_AO22X9 U4958 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ), .D(
        n7282), .Z(n6486) );
  HS65_LL_NAND2X5 U4959 ( .A(n9209), .B(n7120), .Z(n7798) );
  HS65_LL_NAND3X2 U4960 ( .A(n3261), .B(n6125), .C(n8514), .Z(n3262) );
  HS65_LH_NOR2X6 U4961 ( .A(n3233), .B(n8510), .Z(n3234) );
  HS65_LH_IVX9 U4962 ( .A(n8505), .Z(n3228) );
  HS65_LH_NAND3X3 U4963 ( .A(n8535), .B(n8566), .C(n8534), .Z(n8536) );
  HS65_LHS_XNOR2X3 U4964 ( .A(n5913), .B(n5912), .Z(\u_DataPath/toPC2_i [23])
         );
  HS65_LH_NAND2X7 U4965 ( .A(n7678), .B(n7677), .Z(n7754) );
  HS65_LL_AOI12X4 U4966 ( .A(n5910), .B(n5912), .C(n5738), .Z(n5770) );
  HS65_LH_NAND2X7 U4968 ( .A(n3152), .B(n2874), .Z(n8556) );
  HS65_LH_NAND2X7 U4970 ( .A(n3143), .B(n2874), .Z(n8552) );
  HS65_LH_NAND2AX7 U4971 ( .A(n8567), .B(n8568), .Z(n4210) );
  HS65_LL_NOR2X3 U4972 ( .A(n8854), .B(n3403), .Z(n3187) );
  HS65_LL_NOR2X6 U4973 ( .A(n8235), .B(n7921), .Z(n8482) );
  HS65_LH_BFX18 U4974 ( .A(n8288), .Z(n7898) );
  HS65_LH_NOR2X5 U4975 ( .A(n8722), .B(n4712), .Z(n8567) );
  HS65_LL_OAI12X3 U4978 ( .A(n5824), .B(n5827), .C(n5826), .Z(n5912) );
  HS65_LL_NOR2X5 U4979 ( .A(n7797), .B(n7796), .Z(n7120) );
  HS65_LH_NAND2X4 U4980 ( .A(n8044), .B(n8035), .Z(opcode_i[4]) );
  HS65_LH_NAND2X7 U4981 ( .A(n4207), .B(n2866), .Z(n8568) );
  HS65_LH_NOR2X5 U4983 ( .A(n8316), .B(n7868), .Z(n8555) );
  HS65_LHS_XOR2X3 U4984 ( .A(n7753), .B(n7752), .Z(\u_DataPath/pc_4_i [12]) );
  HS65_LHS_XOR2X3 U4985 ( .A(n5774), .B(n5773), .Z(\u_DataPath/toPC2_i [12])
         );
  HS65_LL_NOR2X5 U4987 ( .A(n8049), .B(n8117), .Z(n8635) );
  HS65_LH_NAND2X5 U4988 ( .A(n4714), .B(n8512), .Z(n3233) );
  HS65_LL_NOR3X2 U4989 ( .A(n3413), .B(n8394), .C(n7868), .Z(n3315) );
  HS65_LH_IVX9 U4990 ( .A(n8509), .Z(n3244) );
  HS65_LH_NAND2X5 U4991 ( .A(n7884), .B(\u_DataPath/u_execute/resAdd1_i [16]), 
        .Z(n7865) );
  HS65_LH_NOR2X5 U4992 ( .A(n8835), .B(n4712), .Z(n8497) );
  HS65_LL_AOI12X2 U4993 ( .A(n8119), .B(n8118), .C(n8117), .Z(n8128) );
  HS65_LH_NOR2X6 U4994 ( .A(n8266), .B(n7868), .Z(n8501) );
  HS65_LH_CNIVX3 U4995 ( .A(n4654), .Z(n8495) );
  HS65_LHS_XOR2X3 U4996 ( .A(n6008), .B(n6007), .Z(
        \u_DataPath/u_execute/resAdd1_i [12]) );
  HS65_LH_NOR2X6 U4997 ( .A(\u_DataPath/dataOut_exe_i [27]), .B(n8390), .Z(
        n8558) );
  HS65_LH_NOR2X5 U4998 ( .A(n8387), .B(n9401), .Z(n8531) );
  HS65_LH_NOR2X6 U5000 ( .A(\u_DataPath/dataOut_exe_i [20]), .B(n8390), .Z(
        n8538) );
  HS65_LH_NAND2X4 U5001 ( .A(n4213), .B(n3407), .Z(n3075) );
  HS65_LH_IVX18 U5002 ( .A(\u_DataPath/u_fetch/pc1/N3 ), .Z(n8483) );
  HS65_LH_NAND2X7 U5003 ( .A(n3170), .B(n7869), .Z(n8546) );
  HS65_LL_NOR2AX3 U5006 ( .A(n3055), .B(n3054), .Z(n3056) );
  HS65_LH_NAND2X2 U5007 ( .A(n9376), .B(n8572), .Z(n4188) );
  HS65_LL_AOI12X4 U5008 ( .A(n5902), .B(n5904), .C(n5737), .Z(n5827) );
  HS65_LH_NAND2X7 U5009 ( .A(n3232), .B(n7869), .Z(n8512) );
  HS65_LL_NAND2X2 U5010 ( .A(n9376), .B(n8492), .Z(n3313) );
  HS65_LL_OA12X9 U5011 ( .A(n2932), .B(n3045), .C(n3333), .Z(n3082) );
  HS65_LH_NAND2X4 U5012 ( .A(n3321), .B(n7802), .Z(n8499) );
  HS65_LL_NOR2X5 U5014 ( .A(n7653), .B(n7650), .Z(n7661) );
  HS65_LH_NAND2X7 U5018 ( .A(n6013), .B(n6016), .Z(n5939) );
  HS65_LH_IVX18 U5019 ( .A(n4829), .Z(n7631) );
  HS65_LH_IVX4 U5020 ( .A(n5167), .Z(n7710) );
  HS65_LH_NAND2X7 U5021 ( .A(n5805), .B(n5808), .Z(n5736) );
  HS65_LLS_XOR2X3 U5022 ( .A(n8969), .B(n7089), .Z(n3057) );
  HS65_LH_IVX7 U5023 ( .A(n5716), .Z(n3062) );
  HS65_LL_NOR2X3 U5024 ( .A(n6350), .B(n6342), .Z(n6683) );
  HS65_LL_NOR2X5 U5025 ( .A(n2886), .B(n6149), .Z(n6619) );
  HS65_LH_IVX7 U5026 ( .A(n7905), .Z(n7837) );
  HS65_LL_NOR2X5 U5027 ( .A(n4287), .B(n4286), .Z(n5167) );
  HS65_LL_OAI21X3 U5028 ( .A(n5926), .B(n6034), .C(n5925), .Z(n5962) );
  HS65_LL_NAND2X5 U5029 ( .A(n9111), .B(n3052), .Z(n8262) );
  HS65_LL_OAI21X3 U5030 ( .A(n5724), .B(n5832), .C(n5723), .Z(n5758) );
  HS65_LL_NOR2X6 U5031 ( .A(n6349), .B(n6341), .Z(n6682) );
  HS65_LL_NOR2X5 U5033 ( .A(n6348), .B(n6342), .Z(n6752) );
  HS65_LL_NOR2X5 U5034 ( .A(n6150), .B(n6132), .Z(n6626) );
  HS65_LH_NAND2X4 U5035 ( .A(n5959), .B(n5958), .Z(n5970) );
  HS65_LL_NOR2X5 U5036 ( .A(n6148), .B(n6132), .Z(n6625) );
  HS65_LH_NAND2X5 U5037 ( .A(n5924), .B(n6036), .Z(n5926) );
  HS65_LL_NOR2X3 U5039 ( .A(n8961), .B(n2959), .Z(n2938) );
  HS65_LL_NOR2X5 U5041 ( .A(n2886), .B(n6152), .Z(n6382) );
  HS65_LH_NOR2X5 U5043 ( .A(n8480), .B(n8383), .Z(n8586) );
  HS65_LH_NAND2X4 U5044 ( .A(n5885), .B(n5831), .Z(n5835) );
  HS65_LL_NOR2X6 U5045 ( .A(n2885), .B(n6139), .Z(n6636) );
  HS65_LL_NAND2X2 U5048 ( .A(addr_to_iram[16]), .B(n8692), .Z(n7657) );
  HS65_LH_NAND2X5 U5049 ( .A(n2733), .B(n8391), .Z(n8415) );
  HS65_LH_NAND2X4 U5051 ( .A(n6063), .B(n6062), .Z(n6068) );
  HS65_LH_NAND2X7 U5052 ( .A(addr_to_iram[10]), .B(n8698), .Z(n7647) );
  HS65_LH_NAND2X4 U5053 ( .A(n2733), .B(n8488), .Z(n8444) );
  HS65_LH_NAND2X5 U5054 ( .A(n2733), .B(n8387), .Z(n8457) );
  HS65_LH_NAND2X4 U5055 ( .A(n5819), .B(n5818), .Z(n5823) );
  HS65_LH_IVX7 U5056 ( .A(n2937), .Z(n3041) );
  HS65_LH_NAND2AX4 U5058 ( .A(n8480), .B(n4175), .Z(n7840) );
  HS65_LH_CNIVX3 U5059 ( .A(n8136), .Z(\u_DataPath/cw_memwb_i [0]) );
  HS65_LH_CNIVX3 U5060 ( .A(n8111), .Z(\u_DataPath/cw_tomem_i [8]) );
  HS65_LH_CNIVX3 U5061 ( .A(n8112), .Z(\u_DataPath/cw_tomem_i [7]) );
  HS65_LH_CNIVX3 U5062 ( .A(n8110), .Z(\u_DataPath/cw_tomem_i [6]) );
  HS65_LH_CNIVX3 U5063 ( .A(n8481), .Z(\u_DataPath/cw_tomem_i [0]) );
  HS65_LH_CNIVX3 U5064 ( .A(n8233), .Z(\u_DataPath/jump_i ) );
  HS65_LH_IVX9 U5065 ( .A(n6054), .Z(n5944) );
  HS65_LH_NAND2X7 U5066 ( .A(\u_DataPath/jaddr_i [22]), .B(n8163), .Z(n2885)
         );
  HS65_LH_NAND2X7 U5067 ( .A(n3021), .B(n3404), .Z(n3022) );
  HS65_LH_CNIVX3 U5068 ( .A(n8218), .Z(\u_DataPath/pc_4_to_ex_i [11]) );
  HS65_LH_CNIVX3 U5069 ( .A(n8221), .Z(\u_DataPath/pc_4_to_ex_i [9]) );
  HS65_LH_NAND3X5 U5070 ( .A(n2947), .B(n3030), .C(n8139), .Z(n2949) );
  HS65_LH_CNIVX3 U5071 ( .A(n8216), .Z(\u_DataPath/pc_4_to_ex_i [12]) );
  HS65_LH_CNIVX3 U5072 ( .A(n8222), .Z(\u_DataPath/pc_4_to_ex_i [8]) );
  HS65_LH_CNIVX3 U5073 ( .A(n8214), .Z(\u_DataPath/pc_4_to_ex_i [13]) );
  HS65_LL_NAND4ABX3 U5074 ( .A(n8766), .B(n8763), .C(n2936), .D(n8107), .Z(
        n2937) );
  HS65_LH_CNIVX3 U5075 ( .A(n8223), .Z(\u_DataPath/pc_4_to_ex_i [7]) );
  HS65_LH_CNIVX3 U5076 ( .A(n8213), .Z(\u_DataPath/pc_4_to_ex_i [14]) );
  HS65_LH_CNIVX3 U5077 ( .A(n8224), .Z(\u_DataPath/pc_4_to_ex_i [6]) );
  HS65_LH_CNIVX3 U5078 ( .A(n8212), .Z(\u_DataPath/pc_4_to_ex_i [15]) );
  HS65_LH_CNIVX3 U5079 ( .A(n8225), .Z(\u_DataPath/pc_4_to_ex_i [5]) );
  HS65_LH_CNIVX3 U5080 ( .A(n8211), .Z(\u_DataPath/pc_4_to_ex_i [16]) );
  HS65_LH_CNIVX3 U5081 ( .A(n8209), .Z(\u_DataPath/pc_4_to_ex_i [17]) );
  HS65_LH_CNIVX3 U5082 ( .A(n8208), .Z(\u_DataPath/pc_4_to_ex_i [18]) );
  HS65_LH_CNIVX3 U5083 ( .A(n8226), .Z(\u_DataPath/pc_4_to_ex_i [4]) );
  HS65_LH_CNIVX3 U5084 ( .A(n8206), .Z(\u_DataPath/pc_4_to_ex_i [19]) );
  HS65_LH_CNIVX3 U5085 ( .A(n8205), .Z(\u_DataPath/pc_4_to_ex_i [20]) );
  HS65_LH_CNIVX3 U5086 ( .A(n8204), .Z(\u_DataPath/pc_4_to_ex_i [21]) );
  HS65_LH_CNIVX3 U5087 ( .A(n8227), .Z(\u_DataPath/pc_4_to_ex_i [3]) );
  HS65_LH_NAND2X5 U5088 ( .A(n5859), .B(n5858), .Z(n5861) );
  HS65_LH_CNIVX3 U5089 ( .A(n8219), .Z(\u_DataPath/pc_4_to_ex_i [10]) );
  HS65_LH_CNIVX3 U5090 ( .A(n8202), .Z(\u_DataPath/pc_4_to_ex_i [22]) );
  HS65_LH_CNIVX3 U5091 ( .A(n8229), .Z(\u_DataPath/u_execute/link_value_i [1])
         );
  HS65_LH_CNIVX3 U5093 ( .A(n8200), .Z(\u_DataPath/pc_4_to_ex_i [23]) );
  HS65_LH_CNIVX3 U5094 ( .A(n8198), .Z(\u_DataPath/pc_4_to_ex_i [24]) );
  HS65_LH_CNIVX3 U5095 ( .A(n8197), .Z(\u_DataPath/pc_4_to_ex_i [25]) );
  HS65_LH_CNIVX3 U5097 ( .A(n8196), .Z(\u_DataPath/pc_4_to_ex_i [26]) );
  HS65_LH_CNIVX3 U5098 ( .A(n8194), .Z(\u_DataPath/pc_4_to_ex_i [27]) );
  HS65_LL_NAND2X7 U5099 ( .A(n3030), .B(n8139), .Z(n7618) );
  HS65_LH_CNIVX3 U5100 ( .A(n8193), .Z(\u_DataPath/pc_4_to_ex_i [28]) );
  HS65_LH_CNIVX3 U5101 ( .A(n8191), .Z(\u_DataPath/pc_4_to_ex_i [29]) );
  HS65_LH_CNIVX3 U5102 ( .A(n8190), .Z(\u_DataPath/pc_4_to_ex_i [30]) );
  HS65_LH_CNIVX3 U5103 ( .A(n8289), .Z(\u_DataPath/pc_4_to_ex_i [31]) );
  HS65_LH_IVX44 U5105 ( .A(n3123), .Z(addr_to_iram[12]) );
  HS65_LH_NOR2X6 U5106 ( .A(n6038), .B(n6041), .Z(n6036) );
  HS65_LH_NOR2X5 U5107 ( .A(n6097), .B(n6102), .Z(n5922) );
  HS65_LH_NOR2X5 U5109 ( .A(n5894), .B(n5899), .Z(n5720) );
  HS65_LH_NOR2X6 U5110 ( .A(n7725), .B(n4001), .Z(n7707) );
  HS65_LH_NOR2X6 U5111 ( .A(n5817), .B(n5820), .Z(n5814) );
  HS65_LH_CNIVX3 U5112 ( .A(n9224), .Z(n7722) );
  HS65_LH_NOR2X6 U5113 ( .A(\u_DataPath/jaddr_i [18]), .B(
        \u_DataPath/jaddr_i [20]), .Z(n6326) );
  HS65_LL_IVX7 U5116 ( .A(\u_DataPath/jaddr_i [17]), .Z(n8153) );
  HS65_LH_IVX4 U5117 ( .A(\u_DataPath/dataOut_exe_i [26]), .Z(n3153) );
  HS65_LH_NAND2X7 U5118 ( .A(n8969), .B(n9216), .Z(n6014) );
  HS65_LH_IVX4 U5119 ( .A(n9205), .Z(n7308) );
  HS65_LH_NOR2X5 U5121 ( .A(n8911), .B(n9208), .Z(n5971) );
  HS65_LH_OR2X9 U5123 ( .A(n8944), .B(n9213), .Z(n6109) );
  HS65_LH_IVX9 U5124 ( .A(n8967), .Z(n2940) );
  HS65_LH_IVX4 U5125 ( .A(\u_DataPath/dataOut_exe_i [30]), .Z(n4208) );
  HS65_LH_IVX9 U5126 ( .A(n8966), .Z(n2950) );
  HS65_LL_NOR2X3 U5127 ( .A(n8761), .B(n8764), .Z(n2936) );
  HS65_LH_NAND2X7 U5128 ( .A(n9037), .B(n9212), .Z(n6047) );
  HS65_LH_IVX4 U5130 ( .A(\u_DataPath/dataOut_exe_i [23]), .Z(n3160) );
  HS65_LH_IVX9 U5131 ( .A(n8766), .Z(n8170) );
  HS65_LH_NAND2X5 U5135 ( .A(n9228), .B(n9230), .Z(n4284) );
  HS65_LH_NAND2X7 U5138 ( .A(n9231), .B(n9229), .Z(n4002) );
  HS65_LHS_XNOR2X3 U5139 ( .A(\u_DataPath/jaddr_i [20]), .B(n8968), .Z(n7102)
         );
  HS65_LH_IVX4 U5140 ( .A(\u_DataPath/dataOut_exe_i [15]), .Z(n3273) );
  HS65_LH_NAND2X4 U5142 ( .A(n9039), .B(n9116), .Z(n5897) );
  HS65_LH_CNIVX3 U5145 ( .A(n9221), .Z(n7717) );
  HS65_LH_NAND2X5 U5146 ( .A(n9035), .B(n9115), .Z(n5850) );
  HS65_LH_IVX4 U5147 ( .A(\u_DataPath/dataOut_exe_i [6]), .Z(n3321) );
  HS65_LH_IVX9 U5148 ( .A(\u_DataPath/dataOut_exe_i [16]), .Z(n3205) );
  HS65_LH_NOR2X5 U5150 ( .A(opcode_i[3]), .B(opcode_i[5]), .Z(n7642) );
  HS65_LH_NAND2X7 U5156 ( .A(n7856), .B(n9074), .Z(
        \u_DataPath/dataOut_exe_i [22]) );
  HS65_LL_IVX2 U5157 ( .A(n5681), .Z(n5165) );
  HS65_LL_IVX4 U5158 ( .A(n5679), .Z(n4834) );
  HS65_LL_OAI12X3 U5159 ( .A(n9189), .B(n9073), .C(n8369), .Z(
        \u_DataPath/dataOut_exe_i [24]) );
  HS65_LL_NAND2X4 U5161 ( .A(n5674), .B(n5673), .Z(n5694) );
  HS65_LL_IVX2 U5163 ( .A(n5699), .Z(n5283) );
  HS65_LL_AO12X4 U5165 ( .A(n5160), .B(n5159), .C(n5158), .Z(n5710) );
  HS65_LL_NAND2X2 U5166 ( .A(n7907), .B(n5699), .Z(n7857) );
  HS65_LL_NAND4ABX3 U5167 ( .A(n4453), .B(n5166), .C(n8471), .D(n8470), .Z(
        n4454) );
  HS65_LL_AOI21X3 U5168 ( .A(n5285), .B(n3746), .C(n3745), .Z(n8459) );
  HS65_LL_AOI21X3 U5169 ( .A(n7631), .B(n3813), .C(n3812), .Z(n8460) );
  HS65_LL_NAND2X2 U5170 ( .A(n7907), .B(n4453), .Z(n7842) );
  HS65_LL_AOI12X4 U5171 ( .A(n5285), .B(n3571), .C(n3570), .Z(n8470) );
  HS65_LL_OAI12X3 U5172 ( .A(n5118), .B(n5117), .C(n5116), .Z(n5160) );
  HS65_LH_NAND2X7 U5173 ( .A(n7907), .B(n5686), .Z(n7850) );
  HS65_LL_NAND2X2 U5174 ( .A(n7907), .B(n5166), .Z(n7844) );
  HS65_LL_NAND2X2 U5175 ( .A(n5268), .B(n5267), .Z(n5282) );
  HS65_LL_NAND2X2 U5177 ( .A(n3811), .B(n3810), .Z(n3812) );
  HS65_LL_NAND2X2 U5178 ( .A(n4228), .B(n4227), .Z(n5602) );
  HS65_LL_NOR2AX3 U5179 ( .A(n4452), .B(n4451), .Z(n8471) );
  HS65_LH_AOI21X6 U5180 ( .A(n7631), .B(n4000), .C(n3999), .Z(n8472) );
  HS65_LL_NAND3X2 U5182 ( .A(n4096), .B(n4095), .C(n4094), .Z(n4097) );
  HS65_LL_NAND2X2 U5183 ( .A(n3507), .B(n3506), .Z(n3508) );
  HS65_LL_NAND2X2 U5184 ( .A(n3946), .B(n3945), .Z(n3947) );
  HS65_LL_AOI21X4 U5185 ( .A(n5285), .B(n4141), .C(n4140), .Z(n8468) );
  HS65_LH_NAND2X7 U5186 ( .A(n5643), .B(n4093), .Z(n4094) );
  HS65_LL_OAI21X2 U5188 ( .A(n4863), .B(n5153), .C(n4862), .Z(n4867) );
  HS65_LH_NAND2X7 U5189 ( .A(n5643), .B(n5266), .Z(n5267) );
  HS65_LL_AOI211X3 U5190 ( .A(n3852), .B(n5285), .C(n3851), .D(n3850), .Z(
        n8476) );
  HS65_LH_NAND2X7 U5191 ( .A(n7631), .B(n4057), .Z(n4098) );
  HS65_LL_NAND2X2 U5192 ( .A(n5157), .B(n5156), .Z(n5158) );
  HS65_LLS_XNOR2X3 U5193 ( .A(n4253), .B(n4252), .Z(n4280) );
  HS65_LL_NOR2AX3 U5194 ( .A(n4487), .B(n4486), .Z(n8466) );
  HS65_LL_NAND2AX4 U5195 ( .A(n4139), .B(n4138), .Z(n4140) );
  HS65_LHS_XNOR2X6 U5197 ( .A(n4092), .B(n4091), .Z(n4093) );
  HS65_LLS_XNOR2X3 U5198 ( .A(n3565), .B(n3564), .Z(n3566) );
  HS65_LH_IVX9 U5199 ( .A(n4312), .Z(n4313) );
  HS65_LHS_XNOR2X6 U5201 ( .A(n5199), .B(n5198), .Z(n5222) );
  HS65_LHS_XNOR2X6 U5202 ( .A(n4326), .B(n4325), .Z(n4327) );
  HS65_LH_NAND2X7 U5203 ( .A(n7631), .B(n3902), .Z(n3948) );
  HS65_LL_NOR3X1 U5204 ( .A(n3795), .B(n3794), .C(n3793), .Z(n3796) );
  HS65_LH_NOR2AX3 U5205 ( .A(n3931), .B(n3930), .Z(n3946) );
  HS65_LH_AOI22X6 U5206 ( .A(n9100), .B(n9368), .C(n9187), .D(n8852), .Z(n8297) );
  HS65_LH_OAI12X3 U5209 ( .A(n5611), .B(n2859), .C(n5609), .Z(n5612) );
  HS65_LH_CNIVX3 U5210 ( .A(n8463), .Z(n4791) );
  HS65_LL_NOR2X2 U5211 ( .A(n5634), .B(n5633), .Z(n5635) );
  HS65_LL_NAND3X2 U5213 ( .A(n3886), .B(n3885), .C(n3884), .Z(n3887) );
  HS65_LL_NOR3X1 U5214 ( .A(n3717), .B(n3716), .C(n3715), .Z(n3729) );
  HS65_LL_NOR3X1 U5215 ( .A(n3542), .B(n3541), .C(n3540), .Z(n3569) );
  HS65_LL_NAND4ABX3 U5216 ( .A(n4653), .B(n4652), .C(n4651), .D(n4650), .Z(
        n8467) );
  HS65_LH_NOR3X4 U5217 ( .A(n4898), .B(n4897), .C(n4896), .Z(n4899) );
  HS65_LL_OAI12X3 U5218 ( .A(n3992), .B(n4929), .C(n3991), .Z(n3993) );
  HS65_LH_IVX9 U5219 ( .A(n4536), .Z(n7838) );
  HS65_LL_NOR3X1 U5220 ( .A(n4076), .B(n4075), .C(n4074), .Z(n4096) );
  HS65_LL_IVX2 U5222 ( .A(n4781), .Z(n5119) );
  HS65_LL_NOR3X1 U5223 ( .A(n3989), .B(n3988), .C(n3987), .Z(n3997) );
  HS65_LL_OAI12X2 U5224 ( .A(n4929), .B(n3941), .C(n3940), .Z(n3942) );
  HS65_LH_NOR2AX3 U5225 ( .A(n4054), .B(n4053), .Z(n4055) );
  HS65_LL_NOR2X2 U5226 ( .A(n4137), .B(n4136), .Z(n4138) );
  HS65_LH_NAND2X4 U5229 ( .A(n3804), .B(n5210), .Z(n3806) );
  HS65_LL_NAND2X2 U5231 ( .A(n5643), .B(n4636), .Z(n4651) );
  HS65_LH_NAND2X2 U5233 ( .A(n5615), .B(n4535), .Z(n4278) );
  HS65_LL_NOR3X1 U5234 ( .A(n3978), .B(n3977), .C(n3976), .Z(n3998) );
  HS65_LH_NAND2X5 U5235 ( .A(n5615), .B(n5614), .Z(n5626) );
  HS65_LH_NAND2AX7 U5236 ( .A(n4880), .B(n4879), .Z(n4881) );
  HS65_LH_OAI21X3 U5238 ( .A(n3539), .B(n5646), .C(n3538), .Z(n3540) );
  HS65_LH_OAI21X3 U5239 ( .A(n3713), .B(n4607), .C(n3712), .Z(n3716) );
  HS65_LL_NOR3X1 U5240 ( .A(n5150), .B(n5149), .C(n5148), .Z(n5151) );
  HS65_LH_NAND2X7 U5242 ( .A(n7631), .B(n4908), .Z(n4909) );
  HS65_LH_NOR2X3 U5243 ( .A(n5152), .B(n4895), .Z(n4896) );
  HS65_LH_NAND2X4 U5244 ( .A(n4424), .B(n2867), .Z(n4377) );
  HS65_LH_NAND2X4 U5245 ( .A(n4919), .B(n4916), .Z(n4921) );
  HS65_LH_NAND2X7 U5248 ( .A(n7631), .B(n3854), .Z(n3890) );
  HS65_LH_NOR3X4 U5249 ( .A(n4760), .B(n4759), .C(n4758), .Z(n4779) );
  HS65_LH_NAND2X5 U5250 ( .A(n4555), .B(n4554), .Z(n4556) );
  HS65_LH_NAND2X5 U5254 ( .A(n5632), .B(n5631), .Z(n5634) );
  HS65_LH_OAI12X3 U5255 ( .A(n5241), .B(n4391), .C(n4390), .Z(n4403) );
  HS65_LH_AOI12X2 U5257 ( .A(n4930), .B(n4928), .C(n4927), .Z(n4933) );
  HS65_LH_NOR2X5 U5258 ( .A(n5621), .B(n5226), .Z(n5227) );
  HS65_LH_NOR2X5 U5260 ( .A(n3427), .B(n5204), .Z(n5205) );
  HS65_LL_NOR3X1 U5261 ( .A(n4458), .B(n5321), .C(n4457), .Z(n4475) );
  HS65_LH_AOI21X2 U5263 ( .A(n3939), .B(n4928), .C(n3938), .Z(n3940) );
  HS65_LH_NAND2X5 U5264 ( .A(n4942), .B(n4164), .Z(n3980) );
  HS65_LL_NAND3X2 U5266 ( .A(n4265), .B(n4262), .C(n4260), .Z(n4535) );
  HS65_LH_NAND2X4 U5267 ( .A(n4417), .B(n5631), .Z(n4411) );
  HS65_LH_OAI12X3 U5268 ( .A(n4670), .B(n4669), .C(n4668), .Z(n4695) );
  HS65_LH_NAND2X4 U5269 ( .A(n3751), .B(n5194), .Z(n3753) );
  HS65_LH_OAI21X3 U5272 ( .A(n5646), .B(n4889), .C(n4888), .Z(n4898) );
  HS65_LH_NOR2X3 U5273 ( .A(n5621), .B(n5240), .Z(n3675) );
  HS65_LH_OAI22X3 U5274 ( .A(n4954), .B(n4579), .C(n5146), .D(n3913), .Z(n4603) );
  HS65_LH_IVX7 U5276 ( .A(n4232), .Z(n4233) );
  HS65_LH_NAND2X7 U5277 ( .A(n2733), .B(\u_DataPath/toPC2_i [31]), .Z(n8234)
         );
  HS65_LH_NOR3X3 U5279 ( .A(n4795), .B(n5249), .C(n4163), .Z(n3537) );
  HS65_LH_NOR2X5 U5280 ( .A(n4293), .B(n4317), .Z(n4295) );
  HS65_LH_OAI21X3 U5281 ( .A(n4767), .B(n5656), .C(n4529), .Z(n4530) );
  HS65_LH_AOI22X3 U5282 ( .A(n5229), .B(n4515), .C(n4951), .D(n4560), .Z(n4152) );
  HS65_LH_IVX7 U5283 ( .A(n4839), .Z(n5200) );
  HS65_LL_NAND2X2 U5284 ( .A(n4385), .B(n4384), .Z(n4386) );
  HS65_LH_NAND2X4 U5285 ( .A(n4887), .B(n4148), .Z(n3965) );
  HS65_LH_NAND2X4 U5287 ( .A(n5131), .B(n4560), .Z(n3961) );
  HS65_LH_NAND3X5 U5288 ( .A(n4031), .B(n4030), .C(n4029), .Z(n4032) );
  HS65_LH_NAND2X4 U5289 ( .A(n5661), .B(n4389), .Z(n4347) );
  HS65_LH_AOI21X2 U5290 ( .A(n5618), .B(n5658), .C(n3973), .Z(n3974) );
  HS65_LH_NAND3X5 U5291 ( .A(n5566), .B(n4723), .C(n4722), .Z(n4732) );
  HS65_LH_OAI12X3 U5294 ( .A(n4307), .B(n4332), .C(n4306), .Z(n4308) );
  HS65_LH_NOR2X3 U5295 ( .A(n5621), .B(n4609), .Z(n3717) );
  HS65_LH_NAND3X5 U5296 ( .A(n3866), .B(n3865), .C(n3864), .Z(n3883) );
  HS65_LH_OAI21X3 U5297 ( .A(n5182), .B(n4117), .C(n3601), .Z(n3606) );
  HS65_LH_AOI12X2 U5298 ( .A(n4417), .B(n5630), .C(n4409), .Z(n4410) );
  HS65_LL_NAND3X3 U5299 ( .A(n3491), .B(n4625), .C(n4632), .Z(n3492) );
  HS65_LH_OAI12X3 U5300 ( .A(n5646), .B(n4353), .C(n4352), .Z(n4354) );
  HS65_LH_NAND2X4 U5301 ( .A(n5661), .B(n5243), .Z(n3647) );
  HS65_LH_IVX9 U5305 ( .A(n3923), .Z(n5243) );
  HS65_LL_AOI12X2 U5306 ( .A(n4806), .B(n5672), .C(n4437), .Z(n4438) );
  HS65_LH_NOR3X4 U5308 ( .A(n5466), .B(n5465), .C(n5464), .Z(n5495) );
  HS65_LH_IVX4 U5309 ( .A(n4262), .Z(n4263) );
  HS65_LH_NAND2X7 U5310 ( .A(n4038), .B(n4041), .Z(n3994) );
  HS65_LL_NAND2X2 U5311 ( .A(n4016), .B(n3362), .Z(n3363) );
  HS65_LH_NAND2X5 U5312 ( .A(n4516), .B(n4344), .Z(n4385) );
  HS65_LH_NAND3X3 U5313 ( .A(n5335), .B(n5313), .C(n5402), .Z(n4673) );
  HS65_LH_IVX7 U5314 ( .A(n4319), .Z(n3504) );
  HS65_LH_IVX9 U5315 ( .A(n4435), .Z(n5206) );
  HS65_LH_NOR3X3 U5317 ( .A(n5571), .B(n5471), .C(n5470), .Z(n5472) );
  HS65_LH_IVX4 U5319 ( .A(n4868), .Z(n4803) );
  HS65_LH_NAND2AX7 U5320 ( .A(n3473), .B(n3497), .Z(n4427) );
  HS65_LH_NOR2X5 U5321 ( .A(n4954), .B(n4468), .Z(n3857) );
  HS65_LH_OAI12X3 U5322 ( .A(n9352), .B(n3424), .C(n5423), .Z(n3429) );
  HS65_LH_IVX9 U5324 ( .A(n4806), .Z(n4163) );
  HS65_LL_AOI21X2 U5326 ( .A(n3804), .B(n5211), .C(n3803), .Z(n3805) );
  HS65_LH_NOR2X5 U5327 ( .A(n5287), .B(n5342), .Z(n5352) );
  HS65_LH_NAND2X4 U5328 ( .A(n4942), .B(n4344), .Z(n4058) );
  HS65_LH_NAND2X5 U5329 ( .A(n5131), .B(n4132), .Z(n4133) );
  HS65_LL_NAND2X2 U5330 ( .A(n4040), .B(n3480), .Z(n3475) );
  HS65_LH_NAND2X7 U5331 ( .A(n4303), .B(n4304), .Z(n4232) );
  HS65_LH_NAND2X7 U5332 ( .A(n4259), .B(n4258), .Z(n4950) );
  HS65_LH_OAI21X3 U5333 ( .A(n4939), .B(n4894), .C(n4893), .Z(n4897) );
  HS65_LH_NAND2AX7 U5334 ( .A(n4217), .B(n4316), .Z(n4291) );
  HS65_LH_NAND2X4 U5335 ( .A(n4528), .B(n4344), .Z(n4346) );
  HS65_LH_NOR2X5 U5336 ( .A(n5176), .B(n4558), .Z(n4559) );
  HS65_LH_OAI12X3 U5337 ( .A(n4078), .B(n4077), .C(n4836), .Z(n4079) );
  HS65_LL_IVX2 U5339 ( .A(n4101), .Z(n4645) );
  HS65_LH_NOR2X6 U5341 ( .A(n4077), .B(n4078), .Z(n4391) );
  HS65_LH_OAI12X3 U5343 ( .A(n3800), .B(n3686), .C(n3802), .Z(n3687) );
  HS65_LH_NOR3X4 U5345 ( .A(n5186), .B(n5185), .C(n5184), .Z(n5187) );
  HS65_LH_NOR3X4 U5346 ( .A(n4747), .B(n4746), .C(n4745), .Z(n4780) );
  HS65_LH_AOI22X3 U5347 ( .A(n5234), .B(n4592), .C(n4951), .D(n4617), .Z(n4601) );
  HS65_LH_NAND2X7 U5349 ( .A(n4318), .B(n3471), .Z(n3509) );
  HS65_LH_IVX9 U5350 ( .A(n3872), .Z(n5177) );
  HS65_LH_OAI12X3 U5351 ( .A(n4913), .B(n3895), .C(n4915), .Z(n3896) );
  HS65_LH_IVX9 U5352 ( .A(n3555), .Z(n4873) );
  HS65_LH_AOI21X2 U5354 ( .A(n4490), .B(n5672), .C(n5649), .Z(n3655) );
  HS65_LH_OAI211X5 U5356 ( .A(n4671), .B(n4582), .C(n4129), .D(n4128), .Z(
        n4868) );
  HS65_LL_NAND3X3 U5357 ( .A(n3441), .B(n3440), .C(n4340), .Z(n3872) );
  HS65_LH_NAND2X5 U5358 ( .A(n3910), .B(n3909), .Z(n3911) );
  HS65_LH_NOR2X3 U5359 ( .A(n5603), .B(n3734), .Z(n3737) );
  HS65_LH_OAI12X2 U5360 ( .A(n5603), .B(n3735), .C(n5605), .Z(n3736) );
  HS65_LH_NOR3X4 U5361 ( .A(n3596), .B(n3908), .C(n3595), .Z(n4355) );
  HS65_LH_NAND2X5 U5362 ( .A(n5229), .B(n5170), .Z(n5171) );
  HS65_LH_NOR2X3 U5364 ( .A(n4314), .B(n4318), .Z(n4217) );
  HS65_LH_OAI12X3 U5367 ( .A(n4596), .B(n2897), .C(n4595), .Z(n4597) );
  HS65_LH_NOR2X6 U5368 ( .A(n4064), .B(n4063), .Z(n4113) );
  HS65_LH_NOR2X6 U5369 ( .A(n3460), .B(n3459), .Z(n4849) );
  HS65_LH_NAND2X7 U5371 ( .A(n2733), .B(\u_DataPath/toPC2_i [29]), .Z(n8238)
         );
  HS65_LL_NAND3X3 U5373 ( .A(n3870), .B(n3959), .C(n3790), .Z(n5660) );
  HS65_LH_NAND3X5 U5374 ( .A(n4753), .B(n4752), .C(n4751), .Z(n4759) );
  HS65_LH_NAND3X3 U5375 ( .A(n4763), .B(n4762), .C(n4761), .Z(n4777) );
  HS65_LH_NAND3X5 U5376 ( .A(n5188), .B(n4767), .C(n4766), .Z(n4776) );
  HS65_LH_OAI21X3 U5377 ( .A(n2843), .B(n5129), .C(n4590), .Z(n4077) );
  HS65_LH_NAND2X7 U5378 ( .A(n4316), .B(n4315), .Z(n4326) );
  HS65_LH_NOR2X5 U5379 ( .A(n5399), .B(n5298), .Z(n5402) );
  HS65_LH_NOR2X5 U5380 ( .A(n4320), .B(n4314), .Z(n4290) );
  HS65_LL_AOI21X2 U5381 ( .A(n4538), .B(n3318), .C(n3317), .Z(n4101) );
  HS65_LH_OAI12X3 U5382 ( .A(n4924), .B(n3937), .C(n4926), .Z(n3938) );
  HS65_LL_NOR2X2 U5383 ( .A(n4034), .B(n3990), .Z(n3480) );
  HS65_LH_NAND2X4 U5384 ( .A(n5229), .B(n4356), .Z(n3604) );
  HS65_LL_OAI21X2 U5385 ( .A(n3376), .B(n5179), .C(n5178), .Z(n4437) );
  HS65_LH_IVX7 U5386 ( .A(n4800), .Z(n4132) );
  HS65_LH_NAND2X5 U5387 ( .A(n3934), .B(n3933), .Z(n3943) );
  HS65_LH_NOR2X6 U5388 ( .A(n4011), .B(n3949), .Z(n3362) );
  HS65_LL_IVX4 U5389 ( .A(n3949), .Z(n4017) );
  HS65_LH_CBI4I1X5 U5390 ( .A(n5499), .B(n5572), .C(n5503), .D(n5569), .Z(
        n5488) );
  HS65_LL_NAND3X3 U5392 ( .A(n3985), .B(n3871), .C(n3760), .Z(n5617) );
  HS65_LL_NOR2X3 U5394 ( .A(n3415), .B(n4134), .Z(n4806) );
  HS65_LL_NAND2X4 U5396 ( .A(n3503), .B(n3804), .Z(n4317) );
  HS65_LH_IVX7 U5397 ( .A(n3920), .Z(n3671) );
  HS65_LH_IVX9 U5398 ( .A(n5257), .Z(n3473) );
  HS65_LH_NAND2X5 U5399 ( .A(n5103), .B(n5400), .Z(n5542) );
  HS65_LH_NOR3X4 U5400 ( .A(n4465), .B(n4464), .C(n4463), .Z(n5135) );
  HS65_LH_NOR2X6 U5401 ( .A(n3646), .B(n3645), .Z(n3923) );
  HS65_LH_NOR2X5 U5402 ( .A(n4690), .B(n4702), .Z(n4708) );
  HS65_LH_NOR2X5 U5405 ( .A(n4796), .B(n4582), .Z(n3669) );
  HS65_LH_AOI211X3 U5406 ( .A(n5234), .B(n4750), .C(n4027), .D(n3826), .Z(
        n3828) );
  HS65_LL_NOR2X2 U5407 ( .A(n3932), .B(n4924), .Z(n3478) );
  HS65_LH_NAND2X7 U5408 ( .A(n2892), .B(n5295), .Z(n4864) );
  HS65_LH_NAND2X5 U5409 ( .A(n4904), .B(n4903), .Z(n4907) );
  HS65_LH_NAND3X3 U5410 ( .A(n5502), .B(n5442), .C(n5582), .Z(n4977) );
  HS65_LH_NAND3X3 U5412 ( .A(n4769), .B(n5141), .C(n4768), .Z(n4770) );
  HS65_LH_NAND2X7 U5413 ( .A(n3474), .B(n3359), .Z(n5400) );
  HS65_LH_NOR2X6 U5414 ( .A(\lte_x_59/B[28] ), .B(n3129), .Z(n4333) );
  HS65_LH_NAND2X4 U5415 ( .A(n5292), .B(n5356), .Z(n4690) );
  HS65_LH_IVX7 U5417 ( .A(n3820), .Z(n3822) );
  HS65_LH_NAND2X7 U5419 ( .A(\lte_x_59/B[28] ), .B(n5423), .Z(n4318) );
  HS65_LH_OA12X9 U5420 ( .A(n5126), .B(n4823), .C(n4824), .Z(n2897) );
  HS65_LH_AOI12X2 U5421 ( .A(n5261), .B(n5260), .C(n5259), .Z(n5262) );
  HS65_LH_NAND2X7 U5423 ( .A(n4229), .B(n5569), .Z(n4242) );
  HS65_LH_NAND2X4 U5424 ( .A(\lte_x_59/B[28] ), .B(n4587), .Z(n3649) );
  HS65_LH_NAND2X5 U5425 ( .A(n4878), .B(n4877), .Z(n4884) );
  HS65_LH_IVX4 U5427 ( .A(n3613), .Z(n3614) );
  HS65_LH_IVX4 U5429 ( .A(n4314), .Z(n4315) );
  HS65_LH_AOI21X2 U5430 ( .A(n4943), .B(n4942), .C(n4941), .Z(n4944) );
  HS65_LH_NOR2X6 U5431 ( .A(n4131), .B(n4130), .Z(n4800) );
  HS65_LH_NAND2X5 U5432 ( .A(n4083), .B(n4082), .Z(n4092) );
  HS65_LH_IVX7 U5433 ( .A(n5300), .Z(n5103) );
  HS65_LH_IVX4 U5434 ( .A(n3572), .Z(n3573) );
  HS65_LL_NAND2X2 U5435 ( .A(n5209), .B(n5208), .Z(n5215) );
  HS65_LH_IVX7 U5436 ( .A(n4040), .Z(n3991) );
  HS65_LL_NOR2X3 U5437 ( .A(n3629), .B(n3747), .Z(n3383) );
  HS65_LH_IVX4 U5439 ( .A(n3594), .Z(n3596) );
  HS65_LH_OAI12X3 U5440 ( .A(n5362), .B(n5364), .C(n5290), .Z(n5585) );
  HS65_LH_OAI22X4 U5441 ( .A(n5130), .B(n3756), .C(n4660), .D(n5129), .Z(n3772) );
  HS65_LH_IVX7 U5442 ( .A(n4049), .Z(n3267) );
  HS65_LH_IVX9 U5444 ( .A(n4117), .Z(n4892) );
  HS65_LH_NAND2X4 U5445 ( .A(n5193), .B(n5192), .Z(n5199) );
  HS65_LH_NAND2X5 U5447 ( .A(n4418), .B(n4417), .Z(n4422) );
  HS65_LH_NAND2X7 U5448 ( .A(n3802), .B(n3801), .Z(n3808) );
  HS65_LH_NAND2X4 U5449 ( .A(n4425), .B(n4424), .Z(n4429) );
  HS65_LH_OAI12X3 U5451 ( .A(n3893), .B(n5530), .C(n5506), .Z(n5473) );
  HS65_LH_NAND2X4 U5455 ( .A(n5192), .B(n5290), .Z(n5366) );
  HS65_LHS_XOR2X6 U5456 ( .A(n5126), .B(n4825), .Z(n4826) );
  HS65_LH_NOR2X3 U5457 ( .A(n5004), .B(n2857), .Z(n3954) );
  HS65_LH_NAND2X4 U5458 ( .A(\lte_x_59/B[14] ), .B(n2864), .Z(n4022) );
  HS65_LH_CNIVX3 U5459 ( .A(n3731), .Z(n3732) );
  HS65_LH_OAI22X3 U5461 ( .A(n4671), .B(n2856), .C(n3756), .D(n2843), .Z(n4023) );
  HS65_LH_NAND2X5 U5462 ( .A(\sub_x_53/A[23] ), .B(n4588), .Z(n3718) );
  HS65_LL_OAI22X3 U5464 ( .A(n3756), .B(n4726), .C(n2840), .D(n4583), .Z(n4943) );
  HS65_LH_NAND2X2 U5465 ( .A(\lte_x_59/B[8] ), .B(n2864), .Z(n3674) );
  HS65_LH_NAND2X5 U5468 ( .A(n2842), .B(n4588), .Z(n4060) );
  HS65_LL_NOR2X2 U5470 ( .A(n7834), .B(n2840), .Z(n3420) );
  HS65_LH_NOR2X6 U5471 ( .A(n5320), .B(n5129), .Z(n4798) );
  HS65_LH_IVX9 U5474 ( .A(n4887), .Z(n5146) );
  HS65_LH_OAI21X3 U5475 ( .A(n3365), .B(n5179), .C(n3825), .Z(n3826) );
  HS65_LH_NOR2X3 U5476 ( .A(n4675), .B(n2856), .Z(n3830) );
  HS65_LH_NAND2X4 U5478 ( .A(n4594), .B(n4593), .Z(n4598) );
  HS65_LH_NOR2X3 U5479 ( .A(n2840), .B(n4193), .Z(n4194) );
  HS65_LH_NAND2X7 U5480 ( .A(\lte_x_59/B[24] ), .B(n4551), .Z(n3837) );
  HS65_LH_NAND2X7 U5481 ( .A(\sub_x_53/A[25] ), .B(n2845), .Z(n3836) );
  HS65_LH_IVX7 U5482 ( .A(n4418), .Z(n4409) );
  HS65_LH_NOR2X6 U5483 ( .A(n4984), .B(n5129), .Z(n3907) );
  HS65_LH_IVX4 U5484 ( .A(n5419), .Z(n4417) );
  HS65_LH_NAND2X4 U5486 ( .A(\lte_x_59/B[16] ), .B(n2864), .Z(n4061) );
  HS65_LH_NAND2X5 U5487 ( .A(\lte_x_59/B[21] ), .B(n4587), .Z(n3821) );
  HS65_LH_NAND2X5 U5488 ( .A(n4595), .B(n4561), .Z(n4562) );
  HS65_LH_IVX9 U5489 ( .A(n4951), .Z(n5176) );
  HS65_LH_IVX9 U5490 ( .A(n4341), .Z(n4490) );
  HS65_LH_NAND2X7 U5491 ( .A(\sub_x_53/A[0] ), .B(n4551), .Z(n5183) );
  HS65_LH_OAI21X3 U5492 ( .A(n2871), .B(n5179), .C(n4890), .Z(n4891) );
  HS65_LH_IVX4 U5493 ( .A(n4757), .Z(n4033) );
  HS65_LH_IVX9 U5495 ( .A(n3846), .Z(n4086) );
  HS65_LH_IVX7 U5500 ( .A(n5272), .Z(n5273) );
  HS65_LH_NAND2X5 U5503 ( .A(\sub_x_53/A[29] ), .B(n4588), .Z(n3545) );
  HS65_LH_IVX7 U5504 ( .A(n5258), .Z(n5259) );
  HS65_LH_NAND2X7 U5505 ( .A(n7866), .B(n9065), .Z(
        \u_DataPath/jump_address_i [16]) );
  HS65_LH_NOR2X5 U5506 ( .A(n5656), .B(n5655), .Z(n5657) );
  HS65_LH_NAND2X5 U5507 ( .A(n4206), .B(n4205), .Z(n4226) );
  HS65_LH_NAND2X4 U5508 ( .A(n5313), .B(n5544), .Z(n5325) );
  HS65_LH_NAND2X5 U5511 ( .A(\sub_x_53/A[25] ), .B(n5425), .Z(n3574) );
  HS65_LH_IVX9 U5512 ( .A(n4143), .Z(n3354) );
  HS65_LH_NAND2X7 U5513 ( .A(n2733), .B(\u_DataPath/toPC2_i [27]), .Z(n8240)
         );
  HS65_LH_NAND2X4 U5515 ( .A(n2840), .B(n7623), .Z(n5449) );
  HS65_LH_NAND2X7 U5517 ( .A(n2860), .B(n4967), .Z(n5290) );
  HS65_LH_OAI12X6 U5518 ( .A(n4719), .B(n4718), .C(\sub_x_53/A[25] ), .Z(n5502) );
  HS65_LH_NOR2X5 U5519 ( .A(n4981), .B(n5180), .Z(n5500) );
  HS65_LH_IVX9 U5522 ( .A(n4905), .Z(n3231) );
  HS65_LH_NAND2X5 U5524 ( .A(\sub_x_53/A[29] ), .B(n5422), .Z(n4316) );
  HS65_LH_NOR2X6 U5526 ( .A(\sub_x_53/A[29] ), .B(n5422), .Z(n4314) );
  HS65_LH_NAND2X4 U5528 ( .A(n5327), .B(n5544), .Z(n4666) );
  HS65_LH_NOR2X6 U5530 ( .A(\sub_x_53/A[30] ), .B(n2873), .Z(n4230) );
  HS65_LH_OAI22X4 U5532 ( .A(n7917), .B(n8404), .C(n7915), .D(n8403), .Z(
        \u_DataPath/data_read_ex_1_i [14]) );
  HS65_LH_OAI22X4 U5533 ( .A(n7917), .B(n8343), .C(n7915), .D(n8342), .Z(
        \u_DataPath/data_read_ex_1_i [13]) );
  HS65_LH_OAI22X4 U5534 ( .A(n7902), .B(n8293), .C(n7899), .D(n8183), .Z(
        \u_DataPath/data_read_ex_2_i [12]) );
  HS65_LH_OAI22X4 U5535 ( .A(n7917), .B(n8362), .C(n7915), .D(n8361), .Z(
        \u_DataPath/data_read_ex_1_i [23]) );
  HS65_LH_OAI22X4 U5536 ( .A(n7902), .B(n8415), .C(n7899), .D(n8171), .Z(
        \u_DataPath/data_read_ex_2_i [5]) );
  HS65_LH_OAI22X4 U5537 ( .A(n7917), .B(n8372), .C(n7915), .D(n8371), .Z(
        \u_DataPath/data_read_ex_1_i [24]) );
  HS65_LH_OAI22X4 U5538 ( .A(n7917), .B(n8353), .C(n7915), .D(n8352), .Z(
        \u_DataPath/data_read_ex_1_i [22]) );
  HS65_LH_OAI22X4 U5539 ( .A(n7902), .B(n8304), .C(n7899), .D(n8180), .Z(
        \u_DataPath/data_read_ex_2_i [7]) );
  HS65_LH_OAI22X4 U5540 ( .A(n7902), .B(n8457), .C(n7901), .D(n8386), .Z(
        \u_DataPath/data_read_ex_2_i [18]) );
  HS65_LH_OAI22X4 U5541 ( .A(n7902), .B(n8326), .C(n7900), .D(n8322), .Z(
        \u_DataPath/data_read_ex_2_i [19]) );
  HS65_LH_OAI22X4 U5542 ( .A(n7917), .B(n8378), .C(n7915), .D(n8377), .Z(
        \u_DataPath/data_read_ex_1_i [27]) );
  HS65_LH_OAI22X4 U5543 ( .A(n7902), .B(n8168), .C(n7899), .D(n8156), .Z(
        \u_DataPath/data_read_ex_2_i [1]) );
  HS65_LH_OAI22X4 U5544 ( .A(n7902), .B(n8362), .C(n7899), .D(n8178), .Z(
        \u_DataPath/data_read_ex_2_i [23]) );
  HS65_LH_OAI22X4 U5545 ( .A(n7917), .B(n8358), .C(n7915), .D(n8357), .Z(
        \u_DataPath/data_read_ex_1_i [16]) );
  HS65_LH_OAI22X4 U5546 ( .A(n7902), .B(n8408), .C(n7899), .D(n8175), .Z(
        \u_DataPath/data_read_ex_2_i [17]) );
  HS65_LH_OAI22X4 U5547 ( .A(n7917), .B(n8367), .C(n7915), .D(n8366), .Z(
        \u_DataPath/data_read_ex_1_i [21]) );
  HS65_LH_OAI22X4 U5548 ( .A(n7902), .B(n8321), .C(n7900), .D(n8315), .Z(
        \u_DataPath/data_read_ex_2_i [26]) );
  HS65_LH_OAI22X4 U5549 ( .A(n7902), .B(n8314), .C(n7899), .D(n8310), .Z(
        \u_DataPath/data_read_ex_2_i [6]) );
  HS65_LH_OAI22X4 U5550 ( .A(n7917), .B(n8397), .C(n7915), .D(n8396), .Z(
        \u_DataPath/data_read_ex_1_i [30]) );
  HS65_LH_OAI22X4 U5551 ( .A(n7902), .B(n8330), .C(n7900), .D(n8327), .Z(
        \u_DataPath/data_read_ex_2_i [25]) );
  HS65_LH_OAI22X4 U5552 ( .A(n7902), .B(n8422), .C(n7899), .D(n8158), .Z(
        \u_DataPath/data_read_ex_2_i [31]) );
  HS65_LH_OAI22X4 U5553 ( .A(n7917), .B(n8348), .C(n7915), .D(n8347), .Z(
        \u_DataPath/data_read_ex_1_i [11]) );
  HS65_LH_OAI22X4 U5554 ( .A(n9272), .B(n9186), .C(n9119), .D(n8753), .Z(
        \u_DataPath/data_read_ex_2_i [10]) );
  HS65_LH_OAI22X4 U5555 ( .A(n7902), .B(n8275), .C(n7899), .D(n8261), .Z(
        \u_DataPath/data_read_ex_2_i [8]) );
  HS65_LH_NOR2X5 U5556 ( .A(n4575), .B(n4570), .Z(n3318) );
  HS65_LH_IVX4 U5557 ( .A(n4477), .Z(n4109) );
  HS65_LH_NAND2X7 U5558 ( .A(\lte_x_59/B[14] ), .B(n3366), .Z(n4915) );
  HS65_LH_NOR2X6 U5559 ( .A(\sub_x_53/A[23] ), .B(n5417), .Z(n3698) );
  HS65_LL_IVX7 U5560 ( .A(n3272), .Z(\lte_x_59/B[15] ) );
  HS65_LL_NOR2X5 U5561 ( .A(\lte_x_59/B[16] ), .B(n4985), .Z(n5530) );
  HS65_LH_NOR2X6 U5562 ( .A(\lte_x_59/B[22] ), .B(n5654), .Z(n5603) );
  HS65_LH_NAND2X5 U5563 ( .A(\sub_x_53/A[23] ), .B(n5417), .Z(n3700) );
  HS65_LH_NAND2X7 U5564 ( .A(n2842), .B(n5376), .Z(n4050) );
  HS65_LH_NOR2X6 U5565 ( .A(n3365), .B(n3521), .Z(n3814) );
  HS65_LH_NOR2X3 U5567 ( .A(n5320), .B(n3756), .Z(n3639) );
  HS65_LH_NAND2X7 U5568 ( .A(\lte_x_59/B[21] ), .B(n5418), .Z(n4373) );
  HS65_LH_NAND2X7 U5569 ( .A(\lte_x_59/B[22] ), .B(n5654), .Z(n5605) );
  HS65_LH_NAND2X7 U5571 ( .A(\lte_x_59/B[6] ), .B(n2865), .Z(n4641) );
  HS65_LH_NAND2X7 U5572 ( .A(\sub_x_53/A[20] ), .B(n3376), .Z(n4418) );
  HS65_LH_NOR2X6 U5573 ( .A(\sub_x_53/A[23] ), .B(n4967), .Z(n3731) );
  HS65_LH_NAND2X7 U5574 ( .A(\sub_x_53/A[23] ), .B(n4967), .Z(n3733) );
  HS65_LH_NAND2X7 U5575 ( .A(n2858), .B(n5398), .Z(n4013) );
  HS65_LH_NAND2X5 U5576 ( .A(n5373), .B(n4682), .Z(n5313) );
  HS65_LH_IVX9 U5577 ( .A(n3788), .Z(n5615) );
  HS65_LH_NAND2X7 U5579 ( .A(n2853), .B(n5567), .Z(n3802) );
  HS65_LH_IVX9 U5580 ( .A(\lte_x_59/B[16] ), .Z(n5022) );
  HS65_LH_NOR2X6 U5582 ( .A(\lte_x_59/B[9] ), .B(n5053), .Z(n4876) );
  HS65_LH_NAND2X7 U5583 ( .A(\lte_x_59/B[14] ), .B(n5061), .Z(n4926) );
  HS65_LH_NAND2X7 U5586 ( .A(n2842), .B(n4674), .Z(n4083) );
  HS65_LH_NAND2X7 U5587 ( .A(\lte_x_59/B[6] ), .B(n4147), .Z(n4628) );
  HS65_LH_NOR2X6 U5588 ( .A(n4674), .B(n2842), .Z(n4081) );
  HS65_LH_NAND2X7 U5589 ( .A(n3521), .B(n5048), .Z(n4084) );
  HS65_LHS_XNOR2X3 U5590 ( .A(n5909), .B(n5908), .Z(\u_DataPath/toPC2_i [27])
         );
  HS65_LL_NOR2X3 U5592 ( .A(\lte_x_59/B[14] ), .B(n5061), .Z(n4924) );
  HS65_LH_NOR2X3 U5593 ( .A(n4726), .B(n4795), .Z(n3648) );
  HS65_LH_NAND2X7 U5594 ( .A(\lte_x_59/B[24] ), .B(n3382), .Z(n5193) );
  HS65_LHS_XNOR2X6 U5595 ( .A(n7308), .B(n7307), .Z(
        \u_DataPath/u_execute/link_value_i [28]) );
  HS65_LH_NOR2X6 U5596 ( .A(\lte_x_59/B[24] ), .B(n5180), .Z(n3616) );
  HS65_LH_NOR2X6 U5597 ( .A(n3521), .B(n5048), .Z(n3846) );
  HS65_LH_NAND2X7 U5598 ( .A(n3521), .B(n3365), .Z(n5405) );
  HS65_LH_NOR2X6 U5599 ( .A(n2858), .B(n4683), .Z(n4034) );
  HS65_LH_OA12X9 U5600 ( .A(n4595), .B(n3488), .C(n4594), .Z(n3489) );
  HS65_LH_NAND2X7 U5601 ( .A(n2858), .B(n4683), .Z(n4036) );
  HS65_LH_NAND2X5 U5602 ( .A(n4431), .B(n4516), .Z(n5182) );
  HS65_LH_IVX7 U5603 ( .A(n3488), .Z(n4593) );
  HS65_LH_NAND2X7 U5604 ( .A(\lte_x_59/B[9] ), .B(n5053), .Z(n4878) );
  HS65_LH_NOR2X5 U5605 ( .A(n4581), .B(n3788), .Z(n4528) );
  HS65_LH_IVX9 U5606 ( .A(n8242), .Z(\u_DataPath/branch_target_i [25]) );
  HS65_LH_NOR2X6 U5607 ( .A(n4105), .B(n4108), .Z(n4625) );
  HS65_LHS_XOR2X3 U5608 ( .A(n5752), .B(n5751), .Z(\u_DataPath/toPC2_i [26])
         );
  HS65_LH_IVX9 U5609 ( .A(\lte_x_59/B[1] ), .Z(n4811) );
  HS65_LH_NAND2X7 U5611 ( .A(\lte_x_59/B[4] ), .B(n3352), .Z(n4481) );
  HS65_LH_IVX9 U5612 ( .A(n5418), .Z(n3377) );
  HS65_LH_NOR2X6 U5613 ( .A(\lte_x_59/B[4] ), .B(n3352), .Z(n4100) );
  HS65_LH_IVX9 U5615 ( .A(n5001), .Z(n2870) );
  HS65_LL_NOR2X5 U5616 ( .A(n2925), .B(n3271), .Z(n3272) );
  HS65_LH_IVX9 U5618 ( .A(n5061), .Z(n3366) );
  HS65_LH_NAND2AX7 U5619 ( .A(n4534), .B(n3426), .Z(n3427) );
  HS65_LL_IVX4 U5620 ( .A(n5152), .Z(n4512) );
  HS65_LL_NOR2X2 U5621 ( .A(\lte_x_59/B[7] ), .B(n5312), .Z(n4637) );
  HS65_LL_NOR2X6 U5622 ( .A(n3177), .B(n3176), .Z(\sub_x_53/A[20] ) );
  HS65_LH_NAND2X7 U5624 ( .A(n2733), .B(\u_DataPath/toPC2_i [25]), .Z(n8242)
         );
  HS65_LH_NAND2X5 U5626 ( .A(\lte_x_59/B[8] ), .B(n5373), .Z(n4882) );
  HS65_LL_OR2X18 U5627 ( .A(n3399), .B(n5136), .Z(n3756) );
  HS65_LH_NOR2X6 U5628 ( .A(\lte_x_59/B[4] ), .B(n5032), .Z(n4108) );
  HS65_LH_IVX9 U5630 ( .A(n5423), .Z(n3129) );
  HS65_LH_NOR2X6 U5631 ( .A(\lte_x_59/B[8] ), .B(n5373), .Z(n4880) );
  HS65_LH_NAND2X7 U5633 ( .A(\lte_x_59/B[3] ), .B(n5089), .Z(n4572) );
  HS65_LH_IVX9 U5634 ( .A(n4838), .Z(n4508) );
  HS65_LH_NAND2X5 U5635 ( .A(\lte_x_59/B[3] ), .B(n5321), .Z(n4594) );
  HS65_LH_NAND2X7 U5636 ( .A(n7834), .B(n4550), .Z(n3788) );
  HS65_LH_NOR2X6 U5640 ( .A(\lte_x_59/B[7] ), .B(n5030), .Z(n4622) );
  HS65_LHS_XNOR2X3 U5641 ( .A(n6116), .B(n6115), .Z(
        \u_DataPath/u_execute/resAdd1_i [26]) );
  HS65_LH_IVX9 U5642 ( .A(\u_DataPath/u_idexreg/N16 ), .Z(n8101) );
  HS65_LH_IVX9 U5643 ( .A(n8253), .Z(\u_DataPath/branch_target_i [14]) );
  HS65_LH_IVX9 U5644 ( .A(n8245), .Z(\u_DataPath/branch_target_i [23]) );
  HS65_LHS_XNOR2X3 U5645 ( .A(n5917), .B(n5916), .Z(\u_DataPath/toPC2_i [25])
         );
  HS65_LL_AOI12X4 U5646 ( .A(n5914), .B(n5916), .C(n5739), .Z(n5751) );
  HS65_LL_NAND2X5 U5647 ( .A(n3148), .B(n3147), .Z(n4976) );
  HS65_LH_IVX9 U5648 ( .A(n9052), .Z(n8104) );
  HS65_LL_NAND2X4 U5649 ( .A(n8710), .B(n7780), .Z(n7784) );
  HS65_LL_NAND2X5 U5653 ( .A(n3145), .B(n3144), .Z(n5180) );
  HS65_LH_OAI22X6 U5654 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [24]), .C(
        n8550), .D(n3409), .Z(n3138) );
  HS65_LH_NOR2X5 U5655 ( .A(n8426), .B(n3409), .Z(n3074) );
  HS65_LL_NAND2X5 U5656 ( .A(n3183), .B(n3182), .Z(n5418) );
  HS65_LL_OAI22X3 U5659 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [11]), .C(
        n8345), .D(n3409), .Z(n3072) );
  HS65_LH_OAI22X6 U5661 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [13]), .C(
        n8339), .D(n3409), .Z(n3249) );
  HS65_LH_IVX9 U5662 ( .A(n5425), .Z(n4997) );
  HS65_LL_IVX9 U5663 ( .A(n5321), .Z(n5089) );
  HS65_LH_AOI22X3 U5665 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][2] ), .D(
        n7171), .Z(n6563) );
  HS65_LH_AO22X9 U5666 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ), .D(
        n6635), .Z(n6566) );
  HS65_LH_AO22X9 U5667 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][13] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ), .Z(n6991)
         );
  HS65_LH_AO22X9 U5668 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ), .Z(n6990)
         );
  HS65_LH_AOI22X3 U5669 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ), .D(
        n7285), .Z(n7132) );
  HS65_LH_AOI22X3 U5670 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][13] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][13] ), .Z(n6984)
         );
  HS65_LH_AOI22X3 U5671 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ), .D(
        n7285), .Z(n6876) );
  HS65_LH_AOI22X3 U5673 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ), .D(
        n2888), .Z(n6931) );
  HS65_LH_AOI22X3 U5674 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ), .Z(n6989)
         );
  HS65_LH_AOI22X3 U5675 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ), .Z(n7008)
         );
  HS65_LH_AOI22X3 U5676 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ), .D(
        n7264), .Z(n6932) );
  HS65_LH_AO22X9 U5677 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ), .Z(n7362)
         );
  HS65_LH_AOI22X3 U5679 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][13] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ), .Z(n6988)
         );
  HS65_LH_AOI22X3 U5680 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ), .D(
        n7171), .Z(n6463) );
  HS65_LH_AOI22X3 U5681 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ), .D(
        n2888), .Z(n6889) );
  HS65_LH_AO22X9 U5682 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ), .Z(n7051)
         );
  HS65_LH_AO22X9 U5683 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ), .B(n7429), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ), .Z(n7368)
         );
  HS65_LH_AO22X9 U5685 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ), .D(
        n7282), .Z(n6878) );
  HS65_LH_AO22X9 U5686 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ), .Z(n7056)
         );
  HS65_LH_AO22X9 U5687 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ), .Z(n6970)
         );
  HS65_LH_AO22X9 U5689 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][24] ), .Z(n7572)
         );
  HS65_LH_AO22X9 U5690 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ), .Z(n6971)
         );
  HS65_LH_AO22X9 U5692 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ), .Z(n6778)
         );
  HS65_LH_AOI22X3 U5693 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ), .D(
        n7171), .Z(n6503) );
  HS65_LH_AO22X9 U5694 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][9] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ), .D(
        n7292), .Z(n7137) );
  HS65_LH_AOI22X3 U5695 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ), .D(n7516), 
        .Z(n7251) );
  HS65_LH_AO22X9 U5696 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ), .D(
        n7282), .Z(n6898) );
  HS65_LH_AO22X9 U5697 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ), .D(
        n7586), .Z(n7000) );
  HS65_LH_AOI22X3 U5698 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ), .D(
        n7171), .Z(n7131) );
  HS65_LH_AOI22X3 U5699 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ), .D(
        n7285), .Z(n6896) );
  HS65_LH_AO22X9 U5700 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ), .Z(n7607)
         );
  HS65_LH_AO22X9 U5701 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ), .D(
        n7586), .Z(n6980) );
  HS65_LH_AOI22X3 U5702 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ), .D(
        n6363), .Z(n6869) );
  HS65_LH_AO22X9 U5703 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][25] ), .Z(n7050)
         );
  HS65_LH_AOI22X3 U5705 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ), .D(
        n7264), .Z(n6890) );
  HS65_LH_AO22X9 U5706 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ), .B(n7580), 
        .C(n7579), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ), .Z(n6953) );
  HS65_LH_AO22X9 U5707 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ), .Z(n7581)
         );
  HS65_LH_AO22X9 U5712 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ), .Z(n6976)
         );
  HS65_LH_AO22X9 U5714 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ), .D(
        n7586), .Z(n7040) );
  HS65_LH_AO22X9 U5716 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ), .Z(n7538)
         );
  HS65_LH_AOI22X3 U5717 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ), .D(
        n2889), .Z(n7498) );
  HS65_LH_AO22X9 U5718 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ), .D(n7266), .Z(n6476) );
  HS65_LH_AOI22X3 U5719 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ), .D(
        n7272), .Z(n6913) );
  HS65_LH_AO22X9 U5720 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ), .B(n7429), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ), .Z(n7185)
         );
  HS65_LH_AOI22X3 U5721 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][28] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][28] ), .D(
        n2888), .Z(n6909) );
  HS65_LH_AO22X9 U5722 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ), .D(n7291), .Z(n6490) );
  HS65_LH_AOI22X3 U5724 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ), .D(
        n7171), .Z(n6483) );
  HS65_LH_AOI22X3 U5726 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ), .D(
        n7285), .Z(n6379) );
  HS65_LH_AOI22X3 U5727 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ), .D(
        n7285), .Z(n6916) );
  HS65_LH_AOI22X3 U5728 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ), .D(
        n7171), .Z(n6378) );
  HS65_LH_AO22X9 U5729 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][23] ), .Z(n7235)
         );
  HS65_LH_AO22X9 U5730 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ), .Z(n7036)
         );
  HS65_LH_AOI22X3 U5732 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ), .Z(n7048)
         );
  HS65_LH_AOI22X3 U5733 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ), .D(
        n2889), .Z(n7520) );
  HS65_LH_AOI22X3 U5734 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][23] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ), .D(n7516), 
        .Z(n7231) );
  HS65_LH_AOI22X3 U5735 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ), .D(n7516), 
        .Z(n7191) );
  HS65_LH_AOI22X3 U5736 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][9] ), .D(
        n6363), .Z(n7125) );
  HS65_LH_AO22X9 U5737 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][29] ), .B(n7429), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ), .Z(n7513)
         );
  HS65_LH_AO22X9 U5738 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ), .Z(n7382)
         );
  HS65_LH_AOI22X3 U5739 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ), .D(
        n7264), .Z(n6910) );
  HS65_LH_AO22X9 U5740 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][31] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ), .Z(n6688)
         );
  HS65_LH_AO22X9 U5741 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][14] ), .Z(n7378)
         );
  HS65_LH_AOI22X3 U5742 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][29] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ), .D(
        n2891), .Z(n7515) );
  HS65_LH_AOI22X3 U5743 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ), .Z(n7044)
         );
  HS65_LH_AOI22X3 U5745 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][28] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ), .D(
        n2891), .Z(n7495) );
  HS65_LH_AO22X9 U5747 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ), .Z(n7011)
         );
  HS65_LH_AO22X9 U5748 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][22] ), .Z(n7010)
         );
  HS65_LH_AO22X9 U5749 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ), .D(
        n7586), .Z(n7020) );
  HS65_LH_AO22X9 U5750 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ), .D(
        n7292), .Z(n6861) );
  HS65_LH_AO22X9 U5752 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][3] ), .D(
        n7284), .Z(n6585) );
  HS65_LH_AOI22X3 U5753 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ), .D(
        n7171), .Z(n6583) );
  HS65_LH_AOI22X3 U5754 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][30] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][30] ), .Z(n7420)
         );
  HS65_LH_AOI22X3 U5756 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ), .D(
        n6942), .Z(n6859) );
  HS65_LH_AO22X9 U5757 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ), .B(n7429), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ), .Z(n6328)
         );
  HS65_LH_AOI22X3 U5758 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][19] ), .Z(n6756)
         );
  HS65_LH_AO22X9 U5759 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][7] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ), .Z(n6730)
         );
  HS65_LH_AO22X9 U5761 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ), .Z(n6710)
         );
  HS65_LH_AOI22X3 U5762 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][20] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ), .D(
        n7272), .Z(n6853) );
  HS65_LH_AO22X9 U5763 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ), .Z(n6762)
         );
  HS65_LH_AO22X9 U5765 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ), .D(
        n7282), .Z(n6661) );
  HS65_LH_AO22X9 U5766 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ), .Z(n6761)
         );
  HS65_LH_AOI22X3 U5767 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][18] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ), .D(
        n7285), .Z(n6659) );
  HS65_LH_AOI22X3 U5768 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][18] ), .D(
        n6172), .Z(n6658) );
  HS65_LH_AOI22X3 U5769 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ), .Z(n6760)
         );
  HS65_LH_AOI22X3 U5770 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ), .Z(n6759)
         );
  HS65_LH_AOI22X3 U5771 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ), .D(
        n7285), .Z(n6856) );
  HS65_LH_AOI22X3 U5772 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ), .D(n6740), 
        .Z(n6329) );
  HS65_LH_AOI22X3 U5773 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ), .D(
        n7171), .Z(n6443) );
  HS65_LH_AO22X9 U5774 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ), .Z(n7402)
         );
  HS65_LH_AOI22X3 U5775 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ), .D(n7516), 
        .Z(n7438) );
  HS65_LH_AOI22X3 U5776 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][9] ), .Z(n7028)
         );
  HS65_LH_AOI22X3 U5777 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ), .D(
        n6670), .Z(n7207) );
  HS65_LH_AOI22X3 U5779 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ), .D(n6740), 
        .Z(n7432) );
  HS65_LH_AOI22X3 U5780 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ), .D(
        n6942), .Z(n6406) );
  HS65_LH_AOI22X3 U5781 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][20] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ), .D(
        n2889), .Z(n7478) );
  HS65_LH_AOI22X3 U5782 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ), .D(
        n7171), .Z(n6543) );
  HS65_LH_AOI22X3 U5783 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ), .Z(n7009)
         );
  HS65_LH_AO22X9 U5784 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][12] ), .D(
        n7282), .Z(n6546) );
  HS65_LH_AOI22X3 U5785 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ), .D(
        n7285), .Z(n6403) );
  HS65_LH_AOI22X3 U5787 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ), .D(
        n2891), .Z(n7390) );
  HS65_LH_AO22X9 U5788 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ), .Z(n7486)
         );
  HS65_LH_AO22X9 U5789 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ), .Z(n6357)
         );
  HS65_LH_AO22X9 U5790 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ), .Z(n6356)
         );
  HS65_LH_AOI22X3 U5791 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ), .Z(n6355)
         );
  HS65_LH_AOI22X3 U5792 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][9] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][9] ), .Z(n7024)
         );
  HS65_LH_AOI22X3 U5793 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ), .Z(n6354)
         );
  HS65_LH_AO22X9 U5794 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ), .B(n7580), 
        .C(n7579), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ), .Z(n7347) );
  HS65_LH_AO22X9 U5795 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ), .Z(n7031)
         );
  HS65_LH_AOI22X3 U5797 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ), .D(n7516), 
        .Z(n7211) );
  HS65_LH_AOI22X3 U5798 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ), .D(n2889), .Z(n7393) );
  HS65_LH_AO22X9 U5799 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ), .Z(n7472)
         );
  HS65_LH_AO22X9 U5800 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][9] ), .Z(n7030)
         );
  HS65_LH_AOI22X3 U5802 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][9] ), .Z(n7029)
         );
  HS65_LH_AO22X9 U5804 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ), .Z(n6741)
         );
  HS65_LH_AO22X9 U5805 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][4] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ), .D(
        n7586), .Z(n7351) );
  HS65_LH_AO22X9 U5806 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ), .Z(n7452)
         );
  HS65_LH_AO22X9 U5808 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ), .D(
        n7586), .Z(n7456) );
  HS65_LH_AO22X9 U5809 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][27] ), .Z(n7466)
         );
  HS65_LH_AOI22X3 U5810 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ), .Z(n7068)
         );
  HS65_LH_AO22X9 U5812 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][11] ), .Z(n7070)
         );
  HS65_LH_AO22X9 U5813 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ), .B(n7600), 
        .C(n7599), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ), .Z(n7071)
         );
  HS65_LH_AOI22X3 U5814 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ), .Z(n7064)
         );
  HS65_LH_AO22X9 U5817 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ), .D(
        n7586), .Z(n7060) );
  HS65_LH_AO22X9 U5818 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ), .D(
        n7586), .Z(n6748) );
  HS65_LH_AOI22X3 U5819 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ), .D(
        n2888), .Z(n6849) );
  HS65_LH_AO22X9 U5820 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][16] ), .Z(n7552)
         );
  HS65_LH_AOI22X3 U5822 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ), .D(
        n7264), .Z(n6850) );
  HS65_LH_NOR2X6 U5823 ( .A(opcode_i[5]), .B(n8046), .Z(n8636) );
  HS65_LL_OAI12X3 U5824 ( .A(n5971), .B(n5974), .C(n5973), .Z(n6115) );
  HS65_LH_NOR2X6 U5825 ( .A(n8794), .B(n9050), .Z(\u_DataPath/cw_exmem_i [3])
         );
  HS65_LH_NOR2X6 U5827 ( .A(n9168), .B(n9049), .Z(\u_DataPath/u_idexreg/N15 )
         );
  HS65_LH_OAI21X3 U5828 ( .A(n8871), .B(n9012), .C(n8767), .Z(n8105) );
  HS65_LH_NOR2X6 U5829 ( .A(n8884), .B(n9051), .Z(n8438) );
  HS65_LL_NAND2X4 U5830 ( .A(n3431), .B(n3430), .Z(n4458) );
  HS65_LH_NOR2X6 U5831 ( .A(n8834), .B(n3341), .Z(n3058) );
  HS65_LH_NOR2X6 U5832 ( .A(n8821), .B(n3341), .Z(n4973) );
  HS65_LH_NOR2X6 U5833 ( .A(n8859), .B(n3341), .Z(n3150) );
  HS65_LH_NAND2X7 U5834 ( .A(n8556), .B(n3155), .Z(n3156) );
  HS65_LH_NOR2X5 U5835 ( .A(n8841), .B(n3403), .Z(n3108) );
  HS65_LH_NOR2X6 U5837 ( .A(n8838), .B(n3341), .Z(n3096) );
  HS65_LL_NAND2X2 U5838 ( .A(n3181), .B(n8543), .Z(n3182) );
  HS65_LH_IVX9 U5839 ( .A(n8545), .Z(n3173) );
  HS65_LH_NOR2X6 U5840 ( .A(n3122), .B(n7754), .Z(n7679) );
  HS65_LL_OAI12X3 U5841 ( .A(n5767), .B(n5770), .C(n5769), .Z(n5916) );
  HS65_LHS_XOR2X3 U5843 ( .A(n5771), .B(n5770), .Z(\u_DataPath/toPC2_i [24])
         );
  HS65_LH_NAND2X7 U5844 ( .A(n2733), .B(\u_DataPath/toPC2_i [23]), .Z(n8245)
         );
  HS65_LH_NAND2X7 U5845 ( .A(n2733), .B(\u_DataPath/toPC2_i [14]), .Z(n8253)
         );
  HS65_LL_NAND2X11 U5846 ( .A(n3303), .B(n3302), .Z(n5088) );
  HS65_LH_NAND2X7 U5847 ( .A(n3234), .B(n8511), .Z(n3235) );
  HS65_LH_NOR2X6 U5848 ( .A(n9400), .B(n3341), .Z(n3269) );
  HS65_LL_IVX9 U5850 ( .A(n3340), .Z(n3270) );
  HS65_LH_NAND2X7 U5851 ( .A(n8577), .B(n8318), .Z(n8300) );
  HS65_LH_IVX9 U5852 ( .A(n7764), .Z(n7755) );
  HS65_LH_NAND2X7 U5853 ( .A(n8038), .B(n8039), .Z(n8068) );
  HS65_LH_AOI31X3 U5855 ( .A(n8086), .B(\u_DataPath/immediate_ext_dec_i [1]), 
        .C(n8635), .D(n8085), .Z(n8087) );
  HS65_LH_IVX9 U5856 ( .A(n8277), .Z(\u_DataPath/branch_target_i [7]) );
  HS65_LH_IVX9 U5857 ( .A(n8260), .Z(\u_DataPath/branch_target_i [9]) );
  HS65_LH_IVX7 U5858 ( .A(n8045), .Z(n8046) );
  HS65_LH_IVX9 U5859 ( .A(n8251), .Z(\u_DataPath/branch_target_i [16]) );
  HS65_LH_IVX9 U5860 ( .A(n8247), .Z(\u_DataPath/branch_target_i [21]) );
  HS65_LH_NAND2AX7 U5861 ( .A(\u_DataPath/data_read_ex_2_i [10]), .B(n2874), 
        .Z(n8508) );
  HS65_LH_NOR2X6 U5862 ( .A(n8393), .B(n3340), .Z(n3343) );
  HS65_LL_NAND2X4 U5863 ( .A(n3286), .B(n2874), .Z(n3287) );
  HS65_LH_NAND2X7 U5864 ( .A(n8040), .B(n8039), .Z(n8069) );
  HS65_LH_IVX7 U5865 ( .A(n8519), .Z(n3280) );
  HS65_LH_OAI21X3 U5867 ( .A(n8125), .B(n8124), .C(n8635), .Z(n8127) );
  HS65_LH_OAI21X3 U5868 ( .A(n8075), .B(n8125), .C(n8635), .Z(n8080) );
  HS65_LH_NOR2X6 U5869 ( .A(n8389), .B(n7868), .Z(n8519) );
  HS65_LH_IVX9 U5870 ( .A(n8188), .Z(n8288) );
  HS65_LH_NAND2X7 U5871 ( .A(n2733), .B(\u_DataPath/toPC2_i [16]), .Z(n8251)
         );
  HS65_LH_NAND2X7 U5872 ( .A(n2733), .B(\u_DataPath/toPC2_i [21]), .Z(n8247)
         );
  HS65_LL_NAND3X13 U5873 ( .A(n3333), .B(n3057), .C(n3056), .Z(n3340) );
  HS65_LL_BFX9 U5875 ( .A(n8483), .Z(n7921) );
  HS65_LHS_XOR2X3 U5876 ( .A(n5828), .B(n5827), .Z(\u_DataPath/toPC2_i [22])
         );
  HS65_LH_NOR2X6 U5877 ( .A(n8037), .B(n8117), .Z(n8039) );
  HS65_LH_NOR2X6 U5878 ( .A(n8041), .B(n8117), .Z(n8045) );
  HS65_LH_NAND2X7 U5879 ( .A(n2733), .B(\u_DataPath/toPC2_i [10]), .Z(n8259)
         );
  HS65_LH_NOR2X6 U5880 ( .A(n8047), .B(n8117), .Z(n8634) );
  HS65_LH_NAND2X7 U5881 ( .A(n2733), .B(\u_DataPath/toPC2_i [9]), .Z(n8260) );
  HS65_LH_NAND2X7 U5882 ( .A(n2733), .B(\u_DataPath/toPC2_i [7]), .Z(n8277) );
  HS65_LH_NOR2X6 U5883 ( .A(n7715), .B(n7714), .Z(n7716) );
  HS65_LH_NOR2X6 U5884 ( .A(n8385), .B(n7868), .Z(n8539) );
  HS65_LH_OAI211X3 U5885 ( .A(n8488), .B(n7868), .C(n8487), .D(n8566), .Z(
        n8489) );
  HS65_LH_NOR2X6 U5886 ( .A(n8345), .B(n7868), .Z(n8510) );
  HS65_LH_NAND2X4 U5888 ( .A(n4714), .B(n8535), .Z(n3190) );
  HS65_LH_NOR2X6 U5889 ( .A(n3241), .B(n7868), .Z(n8507) );
  HS65_LH_IVX9 U5891 ( .A(n7671), .Z(n7677) );
  HS65_LH_NOR2X6 U5892 ( .A(n8339), .B(n7868), .Z(n8516) );
  HS65_LH_NAND2X7 U5893 ( .A(n3127), .B(n7869), .Z(n8562) );
  HS65_LH_IVX9 U5896 ( .A(n5791), .Z(n5773) );
  HS65_LH_NAND2X7 U5897 ( .A(n8566), .B(n7306), .Z(n8456) );
  HS65_LH_NAND2X7 U5898 ( .A(n3140), .B(n7869), .Z(n8553) );
  HS65_LH_NAND2X7 U5899 ( .A(n3153), .B(n7869), .Z(n8557) );
  HS65_LHS_XNOR2X6 U5900 ( .A(n5702), .B(n5701), .Z(n5703) );
  HS65_LH_NOR2X6 U5901 ( .A(n8830), .B(n7869), .Z(n3215) );
  HS65_LH_NAND2X7 U5902 ( .A(n7661), .B(n7660), .Z(n7759) );
  HS65_LHS_XNOR2X3 U5903 ( .A(n7713), .B(n7712), .Z(
        \u_DataPath/u_execute/link_value_i [20]) );
  HS65_LH_NAND2X7 U5904 ( .A(n8267), .B(n7869), .Z(n5692) );
  HS65_LH_NAND2X7 U5905 ( .A(n3201), .B(n7869), .Z(n8530) );
  HS65_LH_NAND2X7 U5906 ( .A(n3225), .B(n3407), .Z(n3080) );
  HS65_LH_NOR2X6 U5907 ( .A(n8863), .B(n7869), .Z(n3226) );
  HS65_LH_NAND2X7 U5908 ( .A(n3205), .B(n3407), .Z(n3094) );
  HS65_LH_AOI12X2 U5909 ( .A(n6081), .B(n6083), .C(n6023), .Z(n6024) );
  HS65_LH_NAND2X7 U5910 ( .A(n3242), .B(n7869), .Z(n8509) );
  HS65_LH_NOR2X6 U5911 ( .A(n8849), .B(n7869), .Z(n3257) );
  HS65_LH_NAND2X4 U5912 ( .A(n4714), .B(n8527), .Z(n3206) );
  HS65_LH_IVX9 U5913 ( .A(n5992), .Z(n6007) );
  HS65_LH_NAND2X7 U5915 ( .A(n3252), .B(n7869), .Z(n8518) );
  HS65_LH_NAND2X7 U5916 ( .A(n3273), .B(n7869), .Z(n8524) );
  HS65_LH_NAND2X7 U5917 ( .A(n3188), .B(n7869), .Z(n8535) );
  HS65_LH_NAND2X7 U5919 ( .A(n3336), .B(n7869), .Z(n8496) );
  HS65_LH_NAND2X7 U5920 ( .A(n2733), .B(\u_DataPath/u_fetch/pc1/N3 ), .Z(n8188) );
  HS65_LH_NOR2X5 U5921 ( .A(n8842), .B(n7869), .Z(n3189) );
  HS65_LH_NAND2X7 U5922 ( .A(n7670), .B(n7749), .Z(n7671) );
  HS65_LH_NAND2X7 U5923 ( .A(n2733), .B(\u_DataPath/toPC2_i [3]), .Z(n8281) );
  HS65_LL_OAI12X3 U5924 ( .A(n2879), .B(n3114), .C(n3113), .Z(n8576) );
  HS65_LH_NAND2X7 U5925 ( .A(n2733), .B(\u_DataPath/toPC2_i [4]), .Z(n8280) );
  HS65_LH_IVX9 U5927 ( .A(n7739), .Z(n8161) );
  HS65_LH_IVX9 U5928 ( .A(n7720), .Z(n7723) );
  HS65_LH_NAND2X5 U5929 ( .A(n3205), .B(n7802), .Z(n8527) );
  HS65_LH_NOR2X6 U5931 ( .A(n3120), .B(n7673), .Z(n7660) );
  HS65_LH_NAND2X7 U5932 ( .A(n3307), .B(n7802), .Z(n8492) );
  HS65_LHS_XOR2X6 U5933 ( .A(n7793), .B(n7792), .Z(
        \u_DataPath/u_execute/link_value_i [12]) );
  HS65_LH_NAND2X7 U5934 ( .A(\u_DataPath/dataOut_exe_i [4]), .B(n7802), .Z(
        n3347) );
  HS65_LHS_XOR2X6 U5935 ( .A(n4005), .B(n4004), .Z(n4006) );
  HS65_LH_IVX9 U5936 ( .A(n5999), .Z(n6083) );
  HS65_LH_NAND3X5 U5937 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n4714), .C(
        n7802), .Z(n3283) );
  HS65_LH_NOR2X3 U5938 ( .A(n8833), .B(n7802), .Z(n3134) );
  HS65_LH_NOR2X6 U5941 ( .A(n7691), .B(n7637), .Z(n7739) );
  HS65_LH_IVX9 U5943 ( .A(n5962), .Z(n6077) );
  HS65_LH_NAND2X7 U5944 ( .A(n7730), .B(n7729), .Z(n7792) );
  HS65_LHS_XNOR2X6 U5946 ( .A(n7727), .B(n7729), .Z(
        \u_DataPath/u_execute/link_value_i [10]) );
  HS65_LH_IVX9 U5947 ( .A(n7903), .Z(n5713) );
  HS65_LH_NAND2X5 U5948 ( .A(n9229), .B(n7781), .Z(n7782) );
  HS65_LH_IVX9 U5949 ( .A(n5758), .Z(n5878) );
  HS65_LHS_XNOR2X6 U5950 ( .A(n5901), .B(n5900), .Z(\u_DataPath/toPC2_i [3])
         );
  HS65_LHS_XNOR2X6 U5951 ( .A(n6096), .B(n6095), .Z(
        \u_DataPath/u_execute/resAdd1_i [4]) );
  HS65_LL_NAND2AX7 U5952 ( .A(n3044), .B(n3043), .Z(n3333) );
  HS65_LL_NOR3X4 U5953 ( .A(n2984), .B(n9113), .C(n7640), .Z(n2879) );
  HS65_LH_IVX18 U5954 ( .A(n5234), .Z(n5656) );
  HS65_LL_NOR2X5 U5955 ( .A(n2964), .B(n8262), .Z(n3131) );
  HS65_LL_AOI31X4 U5956 ( .A(n2965), .B(n2961), .C(n2912), .D(n2964), .Z(n3216) );
  HS65_LH_IVX9 U5958 ( .A(n7905), .Z(n7904) );
  HS65_LH_NAND3X5 U5960 ( .A(n2846), .B(n9031), .C(n2946), .Z(n3010) );
  HS65_LH_IVX18 U5961 ( .A(n7906), .Z(n7903) );
  HS65_LH_NAND2X4 U5964 ( .A(n9111), .B(n7085), .Z(n7094) );
  HS65_LH_NOR2X6 U5965 ( .A(n7694), .B(n7775), .Z(n7691) );
  HS65_LH_IVX9 U5966 ( .A(n7690), .Z(n7777) );
  HS65_LH_NAND2X7 U5968 ( .A(n2733), .B(n7854), .Z(n8408) );
  HS65_LH_NOR2X6 U5969 ( .A(n7652), .B(n7647), .Z(n7670) );
  HS65_LL_NOR2X5 U5971 ( .A(n3450), .B(n3449), .Z(n5234) );
  HS65_LH_NAND2X7 U5972 ( .A(n2733), .B(n8345), .Z(n8348) );
  HS65_LH_NOR2X6 U5973 ( .A(n5995), .B(n5998), .Z(n6016) );
  HS65_LL_NOR2X5 U5974 ( .A(n6150), .B(n6140), .Z(n6637) );
  HS65_LL_NAND2X7 U5975 ( .A(n7114), .B(n7113), .Z(n7614) );
  HS65_LH_NAND2X7 U5976 ( .A(n8269), .B(n2980), .Z(n3111) );
  HS65_LH_IVX9 U5979 ( .A(n3314), .Z(n3413) );
  HS65_LH_NOR2X6 U5980 ( .A(n7718), .B(n7787), .Z(n7781) );
  HS65_LL_NOR3X4 U5981 ( .A(n3042), .B(n3041), .C(n3040), .Z(n3043) );
  HS65_LH_IVX7 U5983 ( .A(n3048), .Z(n3049) );
  HS65_LH_BFX18 U5984 ( .A(n8282), .Z(n7882) );
  HS65_LH_NAND2X7 U5985 ( .A(n5930), .B(n5961), .Z(n5932) );
  HS65_LL_NAND2X4 U5987 ( .A(n4713), .B(n9037), .Z(n3395) );
  HS65_LH_NAND2X2 U5988 ( .A(n4713), .B(n9343), .Z(n3164) );
  HS65_LH_OR2X9 U5989 ( .A(\u_DataPath/jaddr_i [18]), .B(n2880), .Z(n6341) );
  HS65_LH_NAND2X4 U5990 ( .A(n4717), .B(n9343), .Z(n4209) );
  HS65_LHS_XNOR2X3 U5991 ( .A(\u_DataPath/jaddr_i [20]), .B(n7618), .Z(n7087)
         );
  HS65_LH_IVX9 U5992 ( .A(n8446), .Z(n7907) );
  HS65_LH_IVX7 U5993 ( .A(n5961), .Z(n5967) );
  HS65_LL_NAND3X3 U5994 ( .A(n2935), .B(n2957), .C(n2963), .Z(n2939) );
  HS65_LH_NAND2X7 U5995 ( .A(n4285), .B(n5688), .Z(n4286) );
  HS65_LH_IVX9 U5996 ( .A(n8591), .Z(n7947) );
  HS65_LL_NOR2X2 U5997 ( .A(n2959), .B(n2958), .Z(n2965) );
  HS65_LL_NOR2X5 U5998 ( .A(n6334), .B(n6353), .Z(n6745) );
  HS65_LH_NAND2X7 U6000 ( .A(n5811), .B(n5814), .Z(n5798) );
  HS65_LL_NOR2X5 U6001 ( .A(n6147), .B(n2886), .Z(n6362) );
  HS65_LH_NAND2X7 U6002 ( .A(n5728), .B(n5757), .Z(n5730) );
  HS65_LH_NAND2X7 U6003 ( .A(n5853), .B(n5718), .Z(n5742) );
  HS65_LH_IVX7 U6005 ( .A(n8393), .Z(n3418) );
  HS65_LH_NAND2X7 U6006 ( .A(n5726), .B(n5779), .Z(n5760) );
  HS65_LL_NOR2X5 U6008 ( .A(n6348), .B(n6334), .Z(n6739) );
  HS65_LH_NAND2X4 U6009 ( .A(n4717), .B(n9341), .Z(n3145) );
  HS65_LL_NOR2X5 U6010 ( .A(n6334), .B(n6349), .Z(n6951) );
  HS65_LH_NAND2X5 U6011 ( .A(n5722), .B(n5834), .Z(n5724) );
  HS65_LH_NAND2X7 U6013 ( .A(n2733), .B(n8265), .Z(n8275) );
  HS65_LH_IVX4 U6014 ( .A(n7665), .Z(n7741) );
  HS65_LH_NAND2X7 U6016 ( .A(\u_DataPath/jaddr_i [25]), .B(n6138), .Z(n6140)
         );
  HS65_LL_NOR2X3 U6017 ( .A(n6349), .B(n6352), .Z(n6689) );
  HS65_LH_NAND2X7 U6019 ( .A(n2733), .B(n8426), .Z(n8449) );
  HS65_LH_NAND2X7 U6020 ( .A(n2733), .B(n8380), .Z(n8397) );
  HS65_LH_NAND2X7 U6021 ( .A(n2733), .B(n8385), .Z(n8412) );
  HS65_LH_IVX9 U6022 ( .A(n7776), .Z(n8084) );
  HS65_LH_NAND2X7 U6025 ( .A(n4713), .B(n8913), .Z(n3346) );
  HS65_LH_NAND2X7 U6026 ( .A(n7695), .B(n7773), .Z(n7775) );
  HS65_LH_IVX9 U6027 ( .A(n8446), .Z(n7906) );
  HS65_LH_NAND2X7 U6029 ( .A(addr_to_iram[4]), .B(n8682), .Z(n7680) );
  HS65_LH_NAND2X7 U6032 ( .A(n5928), .B(n5980), .Z(n5964) );
  HS65_LH_NAND2X7 U6033 ( .A(n4717), .B(n9039), .Z(n3303) );
  HS65_LH_NAND2X7 U6035 ( .A(n5936), .B(n6011), .Z(n5998) );
  HS65_LH_NAND2X7 U6036 ( .A(n2733), .B(n8427), .Z(n8330) );
  HS65_LH_NAND2X7 U6037 ( .A(n2733), .B(n8323), .Z(n8326) );
  HS65_LH_IVX7 U6040 ( .A(n8446), .Z(n7905) );
  HS65_LH_NAND2X7 U6041 ( .A(n2733), .B(n8350), .Z(n8353) );
  HS65_LH_IVX9 U6042 ( .A(n8051), .Z(n8067) );
  HS65_LH_IVX9 U6043 ( .A(n8231), .Z(n8282) );
  HS65_LH_NOR2X6 U6044 ( .A(n5957), .B(n5960), .Z(n5930) );
  HS65_LH_NAND2X7 U6045 ( .A(\u_DataPath/jaddr_i [22]), .B(n8163), .Z(n2886)
         );
  HS65_LH_NAND2X7 U6046 ( .A(n5920), .B(n5919), .Z(n5946) );
  HS65_LL_NAND2X7 U6047 ( .A(n8153), .B(n8152), .Z(n6350) );
  HS65_LH_IVX9 U6048 ( .A(n8052), .Z(n8629) );
  HS65_LH_NOR2X6 U6049 ( .A(n5882), .B(n5887), .Z(n5722) );
  HS65_LL_NAND2X7 U6050 ( .A(\u_DataPath/jaddr_i [17]), .B(n8152), .Z(n6349)
         );
  HS65_LH_NOR2X6 U6051 ( .A(n8090), .B(rst), .Z(
        \u_DataPath/immediate_ext_ex_i [2]) );
  HS65_LH_NAND2X7 U6052 ( .A(n8566), .B(n8264), .Z(n8446) );
  HS65_LH_NAND2X7 U6054 ( .A(n7697), .B(n8055), .Z(n7734) );
  HS65_LH_NOR2X6 U6055 ( .A(n8131), .B(rst), .Z(n8621) );
  HS65_LH_NOR2X6 U6056 ( .A(n8157), .B(rst), .Z(
        \u_DataPath/immediate_ext_ex_i [1]) );
  HS65_LH_NOR2X6 U6058 ( .A(opcode_i[5]), .B(n8070), .Z(n7773) );
  HS65_LH_NOR2X5 U6059 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n8177), .Z(
        n3113) );
  HS65_LH_NOR2X6 U6061 ( .A(n6073), .B(n6078), .Z(n5980) );
  HS65_LH_NAND2X7 U6062 ( .A(n8165), .B(n6131), .Z(n6133) );
  HS65_LH_NOR2X6 U6063 ( .A(n6019), .B(n6022), .Z(n6011) );
  HS65_LH_NAND2X7 U6064 ( .A(n9084), .B(n7643), .Z(n7694) );
  HS65_LH_NOR2X6 U6065 ( .A(n8130), .B(rst), .Z(
        \u_DataPath/immediate_ext_ex_i [0]) );
  HS65_LH_NOR2X6 U6066 ( .A(n5976), .B(n5979), .Z(n5928) );
  HS65_LL_NAND2X7 U6067 ( .A(\u_DataPath/jaddr_i [21]), .B(n8164), .Z(n6148)
         );
  HS65_LH_NAND2X7 U6068 ( .A(n2977), .B(n2976), .Z(n2982) );
  HS65_LH_IVX9 U6069 ( .A(n8050), .Z(n8631) );
  HS65_LH_NAND2X7 U6071 ( .A(\u_DataPath/jaddr_i [19]), .B(n6326), .Z(n2878)
         );
  HS65_LH_IVX44 U6072 ( .A(n3125), .Z(addr_to_iram[13]) );
  HS65_LH_IVX9 U6073 ( .A(n8062), .Z(n8623) );
  HS65_LH_IVX9 U6074 ( .A(n8187), .Z(\u_DataPath/u_idexreg/N31 ) );
  HS65_LH_IVX9 U6076 ( .A(n5915), .Z(n5739) );
  HS65_LH_NAND2X7 U6077 ( .A(n7105), .B(n7104), .Z(n7110) );
  HS65_LH_IVX9 U6078 ( .A(n5812), .Z(n5733) );
  HS65_LL_NAND2X2 U6079 ( .A(n3037), .B(n3036), .Z(n3039) );
  HS65_LH_NAND2X7 U6080 ( .A(n7116), .B(n9234), .Z(n8236) );
  HS65_LL_IVX18 U6081 ( .A(n7758), .Z(addr_to_iram[16]) );
  HS65_LH_IVX9 U6082 ( .A(n8186), .Z(\u_DataPath/u_idexreg/N33 ) );
  HS65_LH_NOR2X6 U6083 ( .A(n4002), .B(n7718), .Z(n4003) );
  HS65_LH_IVX9 U6084 ( .A(n8179), .Z(\u_DataPath/immediate_ext_ex_i [7]) );
  HS65_LH_NOR2X6 U6085 ( .A(n4284), .B(n7728), .Z(n5688) );
  HS65_LH_IVX9 U6086 ( .A(n8185), .Z(\u_DataPath/immediate_ext_ex_i [9]) );
  HS65_LH_IVX9 U6088 ( .A(n8182), .Z(\u_DataPath/immediate_ext_ex_i [10]) );
  HS65_LH_IVX9 U6089 ( .A(n5911), .Z(n5738) );
  HS65_LH_IVX9 U6090 ( .A(n5903), .Z(n5737) );
  HS65_LH_NAND2X7 U6091 ( .A(n7100), .B(n7099), .Z(n7112) );
  HS65_LH_NOR2X6 U6092 ( .A(n4283), .B(n5687), .Z(n4285) );
  HS65_LH_NOR2X6 U6093 ( .A(n5874), .B(n5879), .Z(n5779) );
  HS65_LH_IVX9 U6095 ( .A(n5859), .Z(n5741) );
  HS65_LH_NOR2X6 U6096 ( .A(n6061), .B(n6066), .Z(n5936) );
  HS65_LH_IVX44 U6098 ( .A(n7742), .Z(addr_to_iram[4]) );
  HS65_LH_NOR2X6 U6099 ( .A(n8162), .B(rst), .Z(
        \u_DataPath/immediate_ext_ex_i [3]) );
  HS65_LH_NOR2X6 U6100 ( .A(n5775), .B(n5778), .Z(n5726) );
  HS65_LH_IVX9 U6101 ( .A(n6110), .Z(n5940) );
  HS65_LH_NOR2X2 U6102 ( .A(n8170), .B(rst), .Z(
        \u_DataPath/regfile_addr_out_towb_i [1]) );
  HS65_LH_IVX9 U6103 ( .A(n6106), .Z(n5941) );
  HS65_LH_IVX9 U6104 ( .A(n6114), .Z(n5942) );
  HS65_LH_NOR2X6 U6105 ( .A(n5786), .B(n5772), .Z(n5757) );
  HS65_LH_IVX7 U6107 ( .A(n6082), .Z(n6023) );
  HS65_LH_NAND2X7 U6108 ( .A(n5852), .B(n5851), .Z(n5857) );
  HS65_LH_IVX9 U6109 ( .A(n6118), .Z(n5943) );
  HS65_LH_NOR2X6 U6110 ( .A(n8172), .B(rst), .Z(
        \u_DataPath/immediate_ext_ex_i [5]) );
  HS65_LH_IVX44 U6111 ( .A(n7753), .Z(addr_to_iram[10]) );
  HS65_LH_NOR2X6 U6112 ( .A(n5753), .B(n5756), .Z(n5728) );
  HS65_LH_NOR2X5 U6114 ( .A(n8911), .B(n9204), .Z(n5947) );
  HS65_LH_IVX9 U6117 ( .A(\u_DataPath/dataOut_exe_i [31]), .Z(n4187) );
  HS65_LH_NAND2X4 U6119 ( .A(n9037), .B(n9212), .Z(n5848) );
  HS65_LH_OR2X9 U6120 ( .A(n8969), .B(n9216), .Z(n6013) );
  HS65_LH_OR2X9 U6123 ( .A(n8911), .B(n9203), .Z(n6053) );
  HS65_LH_NAND2X7 U6124 ( .A(n8942), .B(n9222), .Z(n6082) );
  HS65_LH_NAND2X7 U6127 ( .A(n9227), .B(n9225), .Z(n7718) );
  HS65_LH_NOR2X6 U6128 ( .A(n9347), .B(rst), .Z(n8066) );
  HS65_LH_NAND2X4 U6129 ( .A(n9033), .B(n9215), .Z(n5896) );
  HS65_LH_IVX9 U6138 ( .A(\u_DataPath/immediate_ext_dec_i [1]), .Z(n8157) );
  HS65_LL_OR2X9 U6144 ( .A(\u_DataPath/jaddr_i [22]), .B(
        \u_DataPath/jaddr_i [21]), .Z(n6153) );
  HS65_LL_NAND2X7 U6146 ( .A(\u_DataPath/jaddr_i [21]), .B(
        \u_DataPath/jaddr_i [22]), .Z(n6150) );
  HS65_LH_IVX9 U6149 ( .A(\u_DataPath/immediate_ext_dec_i [5]), .Z(n8172) );
  HS65_LH_IVX9 U6154 ( .A(\u_DataPath/dataOut_exe_i [22]), .Z(n3170) );
  HS65_LL_NAND2X5 U6155 ( .A(\u_DataPath/jaddr_i [16]), .B(
        \u_DataPath/jaddr_i [17]), .Z(n6348) );
  HS65_LH_IVX7 U6156 ( .A(n9035), .Z(n3284) );
  HS65_LH_NOR2X6 U6157 ( .A(\u_DataPath/jaddr_i [23]), .B(
        \u_DataPath/jaddr_i [24]), .Z(n6145) );
  HS65_LH_IVX9 U6158 ( .A(\u_DataPath/cw_to_ex_i [19]), .Z(n7874) );
  HS65_LH_OR2X9 U6159 ( .A(n9004), .B(n9209), .Z(n6105) );
  HS65_LH_IVX7 U6160 ( .A(n8944), .Z(n3029) );
  HS65_LH_IVX9 U6161 ( .A(\u_DataPath/dataOut_exe_i [2]), .Z(n3296) );
  HS65_LH_IVX9 U6162 ( .A(n9206), .Z(n7795) );
  HS65_LH_IVX9 U6165 ( .A(n9208), .Z(n7799) );
  HS65_LH_IVX9 U6166 ( .A(n8911), .Z(n3031) );
  HS65_LH_OR2X9 U6167 ( .A(n8911), .B(n9207), .Z(n6113) );
  HS65_LH_IVX9 U6168 ( .A(n9210), .Z(n7797) );
  HS65_LH_IVX9 U6169 ( .A(n9216), .Z(n5696) );
  HS65_LH_NOR2X5 U6170 ( .A(n8911), .B(n9206), .Z(n5952) );
  HS65_LH_IVX9 U6171 ( .A(n9217), .Z(n7713) );
  HS65_LH_NAND2X7 U6172 ( .A(n9218), .B(n9220), .Z(n7711) );
  HS65_LH_NAND2X7 U6175 ( .A(n9116), .B(n9215), .Z(n7725) );
  HS65_LH_NOR2X3 U6176 ( .A(n8913), .B(n9219), .Z(n5839) );
  HS65_LH_IVX9 U6177 ( .A(\u_DataPath/immediate_ext_dec_i [3]), .Z(n8162) );
  HS65_LH_NOR2X6 U6178 ( .A(n8910), .B(rst), .Z(n8283) );
  HS65_LH_IVX9 U6180 ( .A(opcode_i[3]), .Z(n8070) );
  HS65_LH_NAND2X7 U6181 ( .A(n8911), .B(n9208), .Z(n5973) );
  HS65_LH_NAND2X7 U6182 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [12]), 
        .Z(n8052) );
  HS65_LH_NAND2X7 U6183 ( .A(n8911), .B(n9207), .Z(n6114) );
  HS65_LH_NAND2X7 U6184 ( .A(n8911), .B(n9206), .Z(n5954) );
  HS65_LH_NAND2X7 U6185 ( .A(n8685), .B(n8684), .Z(n7644) );
  HS65_LH_NAND2X7 U6186 ( .A(n8680), .B(n8678), .Z(n7645) );
  HS65_LH_NAND2X7 U6187 ( .A(n9181), .B(n9226), .Z(n5863) );
  HS65_LH_NAND2X7 U6188 ( .A(n8911), .B(n9205), .Z(n6118) );
  HS65_LH_NOR2X6 U6189 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(
        \u_DataPath/dataOut_exe_i [1]), .Z(n3112) );
  HS65_LH_NAND2X7 U6191 ( .A(n8911), .B(n9204), .Z(n5949) );
  HS65_LH_IVX9 U6192 ( .A(\u_DataPath/dataOut_exe_i [14]), .Z(n3278) );
  HS65_LH_NAND2X7 U6193 ( .A(n9343), .B(n9203), .Z(n5853) );
  HS65_LH_NAND2X7 U6194 ( .A(n8681), .B(n8679), .Z(n7652) );
  HS65_LH_NAND2X7 U6195 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [13]), 
        .Z(n8064) );
  HS65_LH_NAND2X7 U6197 ( .A(n9145), .B(n9224), .Z(n5755) );
  HS65_LH_NAND2X7 U6198 ( .A(n8911), .B(n9203), .Z(n6054) );
  HS65_LH_NAND2X7 U6200 ( .A(n9342), .B(n9204), .Z(n5859) );
  HS65_LH_IVX9 U6201 ( .A(n9235), .Z(n2977) );
  HS65_LH_IVX9 U6204 ( .A(n9082), .Z(n7643) );
  HS65_LH_NAND2X7 U6206 ( .A(n9343), .B(n9205), .Z(n5745) );
  HS65_LH_NAND2X7 U6207 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [14]), 
        .Z(n8062) );
  HS65_LHS_XNOR2X3 U6209 ( .A(\u_DataPath/jaddr_i [24]), .B(n9077), .Z(n7106)
         );
  HS65_LH_NAND2X7 U6211 ( .A(n9342), .B(n9222), .Z(n5867) );
  HS65_LH_IVX9 U6212 ( .A(opcode_i[1]), .Z(n7697) );
  HS65_LH_NAND2X7 U6214 ( .A(n9342), .B(n9206), .Z(n5907) );
  HS65_LHS_XNOR2X3 U6216 ( .A(\u_DataPath/jaddr_i [23]), .B(n8967), .Z(n7107)
         );
  HS65_LH_NAND2X7 U6218 ( .A(n8706), .B(n8708), .Z(n7686) );
  HS65_LH_NAND2X7 U6220 ( .A(n9341), .B(n9207), .Z(n5750) );
  HS65_LH_NAND2X7 U6221 ( .A(n8705), .B(n8697), .Z(n7658) );
  HS65_LHS_XNOR2X3 U6223 ( .A(\u_DataPath/jaddr_i [25]), .B(n8968), .Z(n7105)
         );
  HS65_LH_NAND2X7 U6224 ( .A(n9341), .B(n9208), .Z(n5915) );
  HS65_LH_NAND2X7 U6225 ( .A(n9343), .B(n9220), .Z(n5812) );
  HS65_LH_NAND2X7 U6226 ( .A(n9343), .B(n9209), .Z(n5769) );
  HS65_LH_NAND2X7 U6227 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [15]), 
        .Z(n8159) );
  HS65_LH_NAND2X7 U6229 ( .A(n9341), .B(n9210), .Z(n5911) );
  HS65_LH_IVX9 U6231 ( .A(\u_DataPath/jaddr_i [24]), .Z(n8151) );
  HS65_LH_IVX9 U6232 ( .A(\u_DataPath/dataOut_exe_i [9]), .Z(n3225) );
  HS65_LH_NAND2X7 U6233 ( .A(n9343), .B(n9213), .Z(n5826) );
  HS65_LH_NAND2X7 U6236 ( .A(n9341), .B(n9217), .Z(n5806) );
  HS65_LH_IVX9 U6237 ( .A(n8932), .Z(n7115) );
  HS65_LH_NOR2X6 U6238 ( .A(\u_DataPath/cw_exmem_i [6]), .B(
        \u_DataPath/cw_exmem_i [4]), .Z(n7098) );
  HS65_LH_NAND2X7 U6240 ( .A(n9343), .B(n9216), .Z(n5903) );
  HS65_LH_IVX9 U6241 ( .A(n9084), .Z(n8055) );
  HS65_LH_NOR2X5 U6242 ( .A(n9075), .B(n8960), .Z(n2941) );
  HS65_LL_IVX4 U6243 ( .A(n9075), .Z(n2942) );
  HS65_LH_NAND2X7 U6244 ( .A(n9004), .B(n9209), .Z(n6106) );
  HS65_LH_IVX7 U6245 ( .A(\u_DataPath/from_mem_data_out_i [5]), .Z(n3331) );
  HS65_LH_NAND2X7 U6248 ( .A(n8944), .B(n9213), .Z(n6110) );
  HS65_LH_NAND2X7 U6250 ( .A(n8943), .B(n9210), .Z(n6028) );
  HS65_LL_IVX7 U6251 ( .A(n8960), .Z(n8139) );
  HS65_LH_IVX9 U6253 ( .A(n9068), .Z(n7695) );
  HS65_LH_NAND2X7 U6254 ( .A(n9267), .B(n9228), .Z(n5788) );
  HS65_LH_NAND2X7 U6255 ( .A(n2733), .B(\u_DataPath/immediate_ext_dec_i [11]), 
        .Z(n8050) );
  HS65_LH_IVX9 U6258 ( .A(Data_out_fromRAM[7]), .Z(n8302) );
  HS65_LL_AOI21X2 U6259 ( .A(n7852), .B(n7853), .C(n7862), .Z(
        \u_DataPath/u_exmemreg/N78 ) );
  HS65_LL_NAND3AX6 U6260 ( .A(n5680), .B(\u_DataPath/cw_to_ex_i [19]), .C(
        n4834), .Z(n5164) );
  HS65_LH_OAI12X3 U6261 ( .A(n9190), .B(n9028), .C(n8340), .Z(
        \u_DataPath/dataOut_exe_i [13]) );
  HS65_LL_NAND4ABX6 U6263 ( .A(n4791), .B(n4790), .C(n4789), .D(n4788), .Z(
        n4792) );
  HS65_LL_NAND2X4 U6264 ( .A(n4370), .B(n8469), .Z(n4455) );
  HS65_LL_NAND2AX4 U6267 ( .A(n5282), .B(n5281), .Z(n5699) );
  HS65_LL_NOR2AX3 U6268 ( .A(n4098), .B(n4097), .Z(n8477) );
  HS65_LL_NAND2AX4 U6270 ( .A(n3744), .B(n3743), .Z(n3745) );
  HS65_LH_OAI12X3 U6271 ( .A(n9189), .B(n8853), .C(n8290), .Z(
        \u_DataPath/dataOut_exe_i [12]) );
  HS65_LH_OAI12X3 U6272 ( .A(n9189), .B(n8887), .C(n8413), .Z(
        \u_DataPath/dataOut_exe_i [5]) );
  HS65_LL_AOI22X1 U6278 ( .A(n8947), .B(n9365), .C(n9187), .D(n9090), .Z(n8267) );
  HS65_LH_NAND2X7 U6279 ( .A(n5285), .B(n4423), .Z(n4452) );
  HS65_LH_OAI12X3 U6281 ( .A(n9189), .B(n9058), .C(n8435), .Z(
        \u_DataPath/dataOut_exe_i [4]) );
  HS65_LL_CNIVX3 U6282 ( .A(n8466), .Z(n5680) );
  HS65_LH_NAND2X7 U6283 ( .A(n5643), .B(n3809), .Z(n3810) );
  HS65_LL_NAND3X2 U6286 ( .A(n5210), .B(n3505), .C(n3495), .Z(n3507) );
  HS65_LHS_XNOR2X6 U6287 ( .A(n5265), .B(n5264), .Z(n5266) );
  HS65_LHS_XNOR2X6 U6288 ( .A(n3808), .B(n3807), .Z(n3809) );
  HS65_LLS_XNOR2X3 U6289 ( .A(n3741), .B(n3740), .Z(n3742) );
  HS65_LL_NAND2X4 U6290 ( .A(n3612), .B(n3611), .Z(n3626) );
  HS65_LH_CNIVX3 U6291 ( .A(n8467), .Z(n4789) );
  HS65_LH_OAI12X3 U6292 ( .A(n3690), .B(n2859), .C(n3689), .Z(n3691) );
  HS65_LLS_XOR2X3 U6293 ( .A(n4056), .B(n4055), .Z(n4057) );
  HS65_LH_NOR2AX3 U6294 ( .A(n4879), .B(n4931), .Z(n4932) );
  HS65_LL_OAI21X2 U6296 ( .A(n3391), .B(n5633), .C(n3390), .Z(n3392) );
  HS65_LL_OA112X4 U6299 ( .A(n5152), .B(n4830), .C(n4831), .D(n2926), .Z(n7848) );
  HS65_LL_OAI21X3 U6300 ( .A(n4420), .B(n5633), .C(n4419), .Z(n4421) );
  HS65_LL_NAND2X2 U6301 ( .A(n3563), .B(n3562), .Z(n3564) );
  HS65_LL_NAND3X2 U6302 ( .A(n5115), .B(n5114), .C(n5113), .Z(n5116) );
  HS65_LH_OAI21X3 U6303 ( .A(n3753), .B(n5633), .C(n3752), .Z(n3754) );
  HS65_LL_OAI21X3 U6304 ( .A(n5530), .B(n5633), .C(n2892), .Z(n3516) );
  HS65_LH_NAND2X7 U6305 ( .A(n4882), .B(n4881), .Z(n4883) );
  HS65_LL_OA12X18 U6306 ( .A(n2929), .B(n3815), .C(n2895), .Z(n5633) );
  HS65_LL_AOI12X2 U6307 ( .A(n4309), .B(n5195), .C(n4308), .Z(n4310) );
  HS65_LH_IVX7 U6308 ( .A(n5195), .Z(n5196) );
  HS65_LL_NAND2X2 U6309 ( .A(n5483), .B(n5482), .Z(n5490) );
  HS65_LH_NOR3X4 U6312 ( .A(n3592), .B(n3591), .C(n3590), .Z(n3612) );
  HS65_LH_NOR2X5 U6313 ( .A(n4088), .B(n4087), .Z(n4089) );
  HS65_LH_NAND2X4 U6314 ( .A(n4845), .B(n3617), .Z(n3563) );
  HS65_LH_NOR3X4 U6315 ( .A(n4403), .B(n4402), .C(n4401), .Z(n4404) );
  HS65_LH_AOI21X2 U6316 ( .A(n6123), .B(n6122), .C(n6121), .Z(n8437) );
  HS65_LH_NOR2AX3 U6320 ( .A(n4235), .B(n4234), .Z(n4236) );
  HS65_LL_NOR2X2 U6321 ( .A(n5060), .B(n5059), .Z(n5070) );
  HS65_LH_OAI21X3 U6322 ( .A(n4119), .B(n4855), .C(n3523), .Z(n3542) );
  HS65_LL_NOR3X1 U6323 ( .A(n3883), .B(n3882), .C(n3881), .Z(n3884) );
  HS65_LL_NOR2X2 U6324 ( .A(n5481), .B(n5480), .Z(n5483) );
  HS65_LH_OAI21X3 U6325 ( .A(n5226), .B(n4855), .C(n3914), .Z(n3929) );
  HS65_LH_OAI12X3 U6326 ( .A(n4921), .B(n3815), .C(n4920), .Z(n4922) );
  HS65_LH_NOR2AX3 U6328 ( .A(n4086), .B(n4085), .Z(n4087) );
  HS65_LL_NAND3X3 U6329 ( .A(n4780), .B(n4779), .C(n4778), .Z(n4781) );
  HS65_LH_AOI12X2 U6330 ( .A(n4043), .B(n4879), .C(n4042), .Z(n4044) );
  HS65_LH_NOR2X6 U6331 ( .A(n4844), .B(n4843), .Z(n5153) );
  HS65_LH_NAND2X2 U6333 ( .A(n5285), .B(n5284), .Z(n5597) );
  HS65_LH_OAI21X3 U6334 ( .A(n4744), .B(n5656), .C(n4272), .Z(n4273) );
  HS65_LL_NAND3X2 U6336 ( .A(n3678), .B(n3677), .C(n3676), .Z(n3679) );
  HS65_LH_NAND2X4 U6340 ( .A(n3618), .B(n4879), .Z(n3493) );
  HS65_LL_OA12X4 U6341 ( .A(n3816), .B(n3370), .C(n3369), .Z(n2895) );
  HS65_LH_NAND3X3 U6342 ( .A(n4179), .B(n4178), .C(n4177), .Z(n4204) );
  HS65_LH_AOI21X2 U6343 ( .A(n5234), .B(n4765), .C(n4354), .Z(n4360) );
  HS65_LL_OAI12X2 U6344 ( .A(n5102), .B(n5101), .C(n5100), .Z(n5111) );
  HS65_LH_IVX9 U6345 ( .A(n3589), .Z(n4895) );
  HS65_LH_OAI12X3 U6346 ( .A(n3462), .B(n5621), .C(n3461), .Z(n3463) );
  HS65_LH_NAND2X4 U6348 ( .A(n3426), .B(n4504), .Z(n4607) );
  HS65_LH_OAI21X3 U6350 ( .A(n4954), .B(n3962), .C(n3961), .Z(n3978) );
  HS65_LH_OAI21X3 U6352 ( .A(n4220), .B(n4319), .C(n4219), .Z(n4221) );
  HS65_LH_OAI21X3 U6353 ( .A(n3975), .B(n5656), .C(n3974), .Z(n3976) );
  HS65_LH_NAND3AX6 U6357 ( .A(n5664), .B(n5663), .C(n5662), .Z(n5665) );
  HS65_LH_NAND2X7 U6358 ( .A(n4149), .B(n4162), .Z(n5614) );
  HS65_LH_NOR3X3 U6359 ( .A(n5089), .B(n4458), .C(n4457), .Z(n3845) );
  HS65_LL_OAI12X2 U6361 ( .A(n5018), .B(n5017), .C(n5016), .Z(n5019) );
  HS65_LH_OAI21X3 U6362 ( .A(n5182), .B(n5226), .C(n3647), .Z(n3681) );
  HS65_LH_CNIVX3 U6363 ( .A(n5577), .Z(n5581) );
  HS65_LH_OAI21X3 U6364 ( .A(n4954), .B(n4953), .C(n4952), .Z(n4957) );
  HS65_LH_OAI21X3 U6365 ( .A(n5177), .B(n4842), .C(n4432), .Z(n4433) );
  HS65_LH_NAND2X7 U6369 ( .A(n4051), .B(n4916), .Z(n4052) );
  HS65_LH_NAND2X5 U6370 ( .A(n6123), .B(n4381), .Z(n4135) );
  HS65_LH_NOR2AX3 U6371 ( .A(n4072), .B(n4071), .Z(n4073) );
  HS65_LH_AOI21X2 U6373 ( .A(n4951), .B(n5142), .C(n3859), .Z(n3885) );
  HS65_LH_NAND2AX7 U6374 ( .A(n4121), .B(n4384), .Z(n4388) );
  HS65_LL_NOR2X2 U6375 ( .A(n3375), .B(n4419), .Z(n3381) );
  HS65_LH_IVX9 U6376 ( .A(n8234), .Z(\u_DataPath/branch_target_i [31]) );
  HS65_LH_NAND2X7 U6377 ( .A(n3557), .B(n3556), .Z(n4816) );
  HS65_LH_OAI12X3 U6378 ( .A(n5200), .B(n4842), .C(n4841), .Z(n4843) );
  HS65_LH_NAND3X3 U6379 ( .A(n3917), .B(n3916), .C(n3915), .Z(n3918) );
  HS65_LH_NOR3X3 U6380 ( .A(n4581), .B(n5152), .C(n4025), .Z(n4026) );
  HS65_LH_OAI21X3 U6381 ( .A(n3584), .B(n3101), .C(n3583), .Z(n3591) );
  HS65_LH_CNIVX3 U6382 ( .A(n5486), .Z(n5305) );
  HS65_LH_NAND2X4 U6383 ( .A(n5174), .B(n5229), .Z(n3827) );
  HS65_LH_IVX9 U6384 ( .A(n4025), .Z(n4504) );
  HS65_LH_OAI21X3 U6386 ( .A(n4737), .B(n5656), .C(n4392), .Z(n4402) );
  HS65_LH_NOR2X5 U6387 ( .A(n3762), .B(n3599), .Z(n3600) );
  HS65_LH_NOR3X1 U6388 ( .A(n5476), .B(n5511), .C(n5475), .Z(n5477) );
  HS65_LH_NAND2X4 U6389 ( .A(n4887), .B(n4873), .Z(n4124) );
  HS65_LL_NOR3X1 U6390 ( .A(n4777), .B(n4776), .C(n4775), .Z(n4778) );
  HS65_LH_AOI22X3 U6391 ( .A(n4887), .B(n4839), .C(n4951), .D(n4835), .Z(n3842) );
  HS65_LL_NAND2AX4 U6393 ( .A(n3476), .B(n3475), .Z(n4928) );
  HS65_LH_AOI22X3 U6394 ( .A(n5144), .B(n4616), .C(n4887), .D(n4007), .Z(n4008) );
  HS65_LH_AOI22X3 U6395 ( .A(n5229), .B(n4176), .C(n5618), .D(n4614), .Z(n4009) );
  HS65_LL_AOI22X1 U6396 ( .A(\sub_x_53/A[30] ), .B(n4493), .C(n5672), .D(n4492), .Z(n5704) );
  HS65_LH_IVX9 U6397 ( .A(n4420), .Z(n5631) );
  HS65_LH_OAI21X3 U6398 ( .A(n5653), .B(n5652), .C(n5651), .Z(n5664) );
  HS65_LH_AOI21X2 U6399 ( .A(n5659), .B(n5658), .C(n5657), .Z(n5663) );
  HS65_LH_OAI21X3 U6400 ( .A(n4749), .B(n5656), .C(n4461), .Z(n4471) );
  HS65_LH_NAND2X4 U6401 ( .A(n4951), .B(n5143), .Z(n4466) );
  HS65_LHS_XNOR2X6 U6403 ( .A(n4478), .B(n4632), .Z(n4479) );
  HS65_LHS_XOR2X6 U6404 ( .A(n3853), .B(n3815), .Z(n3854) );
  HS65_LH_AOI21X2 U6405 ( .A(n3505), .B(n5211), .C(n3504), .Z(n3506) );
  HS65_LL_OAI112X1 U6406 ( .A(n4954), .B(n4070), .C(n4069), .D(n4068), .Z(
        n4071) );
  HS65_LH_AOI21X2 U6407 ( .A(n4491), .B(n4508), .C(n4263), .Z(n4264) );
  HS65_LH_OAI21X3 U6408 ( .A(n4740), .B(n5656), .C(n4058), .Z(n4076) );
  HS65_LL_IVX4 U6409 ( .A(n3894), .Z(n4916) );
  HS65_LH_NAND3X3 U6410 ( .A(n5509), .B(n4705), .C(n4704), .Z(n4706) );
  HS65_LL_AOI12X2 U6411 ( .A(n4937), .B(n4887), .C(n2901), .Z(n4555) );
  HS65_LH_OAI21X3 U6412 ( .A(n4439), .B(n4700), .C(n4438), .Z(n4440) );
  HS65_LH_NOR2X6 U6414 ( .A(n3878), .B(n3877), .Z(n5204) );
  HS65_LH_NAND2X5 U6416 ( .A(n5618), .B(n5206), .Z(n4856) );
  HS65_LH_OAI12X3 U6417 ( .A(n4499), .B(n4498), .C(n4836), .Z(n4511) );
  HS65_LH_IVX9 U6418 ( .A(n4614), .Z(n5226) );
  HS65_LH_OAI21X3 U6420 ( .A(n3534), .B(n5656), .C(n3533), .Z(n3541) );
  HS65_LL_NOR2X2 U6421 ( .A(n4992), .B(n4977), .Z(n5115) );
  HS65_LH_OAI21X3 U6422 ( .A(n4117), .B(n4838), .C(n4079), .Z(n4349) );
  HS65_LH_NAND2X4 U6423 ( .A(n4951), .B(n4937), .Z(n3986) );
  HS65_LH_NAND2X5 U6424 ( .A(n4836), .B(n4148), .Z(n4162) );
  HS65_LH_OAI21X3 U6425 ( .A(n5188), .B(n5656), .C(n5187), .Z(n5189) );
  HS65_LH_NAND2X4 U6427 ( .A(n4951), .B(n4950), .Z(n4952) );
  HS65_LH_AOI22X3 U6428 ( .A(n5234), .B(n4764), .C(n5144), .D(n4937), .Z(n4151) );
  HS65_LL_NAND2X4 U6429 ( .A(n4037), .B(n3480), .Z(n3935) );
  HS65_LH_NAND2AX7 U6430 ( .A(n4946), .B(n2898), .Z(n4947) );
  HS65_LH_IVX9 U6431 ( .A(n4919), .Z(n3282) );
  HS65_LL_NAND3X3 U6432 ( .A(n3985), .B(n3984), .C(n3983), .Z(n4937) );
  HS65_LH_NAND2X4 U6433 ( .A(n5659), .B(n4872), .Z(n3583) );
  HS65_LH_AOI21X2 U6434 ( .A(n3737), .B(n5607), .C(n3736), .Z(n3738) );
  HS65_LH_AND2X4 U6436 ( .A(n2733), .B(\u_DataPath/toPC2_i [30]), .Z(
        \u_DataPath/branch_target_i [30]) );
  HS65_LL_NAND2X2 U6437 ( .A(n3875), .B(n3876), .Z(n3402) );
  HS65_LH_IVX9 U6439 ( .A(n4513), .Z(n5658) );
  HS65_LH_NOR2X6 U6440 ( .A(n4255), .B(n4254), .Z(n4955) );
  HS65_LL_NAND2AX4 U6441 ( .A(n3458), .B(n3457), .Z(n5174) );
  HS65_LH_OAI21X3 U6442 ( .A(n5656), .B(n5141), .C(n5140), .Z(n5149) );
  HS65_LL_NAND3X2 U6443 ( .A(n3960), .B(n3959), .C(n3958), .Z(n4560) );
  HS65_LH_NAND2X4 U6444 ( .A(n5661), .B(n5617), .Z(n3761) );
  HS65_LH_NAND2X4 U6448 ( .A(n4516), .B(n4872), .Z(n4080) );
  HS65_LH_NAND2X2 U6449 ( .A(n4887), .B(n4886), .Z(n4888) );
  HS65_LH_OAI12X3 U6451 ( .A(n4681), .B(n4680), .C(n4679), .Z(n4689) );
  HS65_LH_AOI21X2 U6452 ( .A(n5618), .B(n4393), .C(n3532), .Z(n3533) );
  HS65_LH_NAND2X2 U6453 ( .A(n3426), .B(n5660), .Z(n4519) );
  HS65_LH_OAI12X3 U6454 ( .A(n4575), .B(n4574), .C(n4573), .Z(n4576) );
  HS65_LH_AOI21X2 U6455 ( .A(n4017), .B(n4016), .C(n5466), .Z(n4018) );
  HS65_LH_NAND2X4 U6456 ( .A(n5144), .B(n5142), .Z(n4467) );
  HS65_LH_AND2X4 U6457 ( .A(n5234), .B(n3451), .Z(n3452) );
  HS65_LL_AO12X4 U6461 ( .A(n5274), .B(n3374), .C(n3373), .Z(n5630) );
  HS65_LH_AOI21X2 U6462 ( .A(n5582), .B(n5580), .C(n5013), .Z(n5017) );
  HS65_LL_NOR2AX3 U6463 ( .A(n3921), .B(n3671), .Z(n4609) );
  HS65_LH_IVX9 U6464 ( .A(n8238), .Z(\u_DataPath/branch_target_i [29]) );
  HS65_LH_NAND2X5 U6465 ( .A(n3426), .B(n4120), .Z(n4384) );
  HS65_LL_OAI12X2 U6466 ( .A(n5081), .B(n5011), .C(n5010), .Z(n5020) );
  HS65_LH_AOI22X3 U6467 ( .A(n5131), .B(n5142), .C(n4942), .D(n3872), .Z(n3843) );
  HS65_LH_OAI12X3 U6468 ( .A(n3969), .B(n3757), .C(n5672), .Z(n3799) );
  HS65_LH_IVX4 U6469 ( .A(n3876), .Z(n3877) );
  HS65_LH_NAND2X4 U6470 ( .A(n5443), .B(n3630), .Z(n3638) );
  HS65_LL_IVX2 U6471 ( .A(n4014), .Z(n3246) );
  HS65_LH_NAND3X2 U6472 ( .A(n4852), .B(n4851), .C(n5178), .Z(n4853) );
  HS65_LH_NAND2AX7 U6473 ( .A(n3520), .B(n3519), .Z(n4872) );
  HS65_LH_OAI21X2 U6475 ( .A(n2873), .B(n5179), .C(n5178), .Z(n4527) );
  HS65_LL_NOR2X2 U6476 ( .A(n3483), .B(n4629), .Z(n3484) );
  HS65_LL_NOR2X3 U6477 ( .A(n3863), .B(n3862), .Z(n4435) );
  HS65_LL_NAND2X4 U6478 ( .A(n3586), .B(n3585), .Z(n4120) );
  HS65_LH_AOI21X2 U6479 ( .A(n5275), .B(n5274), .C(n5273), .Z(n5276) );
  HS65_LL_NOR2X2 U6481 ( .A(n4257), .B(n4256), .Z(n4953) );
  HS65_LH_OAI12X3 U6482 ( .A(n4015), .B(n4011), .C(n4013), .Z(n3364) );
  HS65_LL_NAND3X3 U6483 ( .A(n4591), .B(n3674), .C(n3673), .Z(n4176) );
  HS65_LL_NAND2X4 U6484 ( .A(n5304), .B(n3893), .Z(n5522) );
  HS65_LH_NAND3X3 U6485 ( .A(n3531), .B(n5178), .C(n3530), .Z(n3532) );
  HS65_LL_NOR3X1 U6486 ( .A(n3434), .B(n3982), .C(n3433), .Z(n5172) );
  HS65_LH_NAND2X7 U6487 ( .A(n5009), .B(n5507), .Z(n5081) );
  HS65_LH_NAND2X4 U6488 ( .A(n5270), .B(n5467), .Z(n5082) );
  HS65_LL_NOR2X2 U6489 ( .A(n4524), .B(n3834), .Z(n3835) );
  HS65_LH_OAI12X3 U6491 ( .A(n4725), .B(n4795), .C(n3759), .Z(n4254) );
  HS65_LH_NAND3X3 U6492 ( .A(n3972), .B(n3971), .C(n3970), .Z(n3973) );
  HS65_LH_OAI21X3 U6494 ( .A(n4197), .B(n4196), .C(n4195), .Z(n4198) );
  HS65_LH_OAI21X3 U6495 ( .A(n4798), .B(n4797), .C(n5131), .Z(n4799) );
  HS65_LH_IVX4 U6497 ( .A(n3841), .Z(n3781) );
  HS65_LH_NAND2X5 U6498 ( .A(n5434), .B(n4408), .Z(n4413) );
  HS65_LH_NAND2X5 U6499 ( .A(n3474), .B(n3359), .Z(n4015) );
  HS65_LH_AOI21X6 U6500 ( .A(\sub_x_53/A[2] ), .B(n2864), .C(n4798), .Z(n3519)
         );
  HS65_LH_NAND2X4 U6502 ( .A(n4143), .B(n4099), .Z(n4104) );
  HS65_LL_OAI12X3 U6503 ( .A(n2892), .B(n3515), .C(n5531), .Z(n5274) );
  HS65_LH_NAND2X4 U6505 ( .A(n4013), .B(n4012), .Z(n4021) );
  HS65_LH_NAND2X4 U6508 ( .A(n3733), .B(n3732), .Z(n3741) );
  HS65_LL_OAI12X2 U6509 ( .A(n5269), .B(n5272), .C(n5270), .Z(n3373) );
  HS65_LH_CBI4I1X5 U6510 ( .A(n4102), .B(n4099), .C(n3354), .D(n3353), .Z(
        n3356) );
  HS65_LH_OAI211X3 U6511 ( .A(n5652), .B(n4582), .C(n3603), .D(n3602), .Z(
        n4356) );
  HS65_LH_NAND2X4 U6512 ( .A(n4915), .B(n4914), .Z(n4923) );
  HS65_LL_AOI12X3 U6513 ( .A(n3497), .B(n5260), .C(n3496), .Z(n4426) );
  HS65_LL_NAND2AX4 U6514 ( .A(n3351), .B(n4638), .Z(n3358) );
  HS65_LH_NOR2X6 U6515 ( .A(n3613), .B(n3616), .Z(n3804) );
  HS65_LH_NAND2X4 U6516 ( .A(n5605), .B(n5604), .Z(n5613) );
  HS65_LH_NAND2X4 U6517 ( .A(n4846), .B(n4845), .Z(n4847) );
  HS65_LH_CNIVX3 U6518 ( .A(n4037), .Z(n3992) );
  HS65_LH_NAND2X4 U6520 ( .A(n3474), .B(n4544), .Z(n3457) );
  HS65_LH_NAND2X2 U6521 ( .A(n4572), .B(n4571), .Z(n4577) );
  HS65_LH_OAI12X3 U6522 ( .A(n4581), .B(n4580), .C(n3529), .Z(n4804) );
  HS65_LH_AOI21X6 U6523 ( .A(\sub_x_53/A[2] ), .B(n4544), .C(n4541), .Z(n3876)
         );
  HS65_LH_CNIVX3 U6524 ( .A(n4927), .Z(n3937) );
  HS65_LH_NAND2X4 U6525 ( .A(n5275), .B(n5271), .Z(n5277) );
  HS65_LH_NAND2X4 U6526 ( .A(n4507), .B(n4516), .Z(n4608) );
  HS65_LH_IVX7 U6527 ( .A(n3491), .Z(n3483) );
  HS65_LH_NAND2X4 U6528 ( .A(n3833), .B(n3984), .Z(n3770) );
  HS65_LH_CNIVX3 U6529 ( .A(n3907), .Z(n3664) );
  HS65_LH_IVX9 U6533 ( .A(n3969), .Z(n4134) );
  HS65_LH_NOR2X3 U6534 ( .A(n4795), .B(n4660), .Z(n3640) );
  HS65_LH_OAI21X3 U6535 ( .A(n4981), .B(n4795), .C(n3603), .Z(n3551) );
  HS65_LH_AOI21X2 U6536 ( .A(\sub_x_53/A[17] ), .B(n4588), .C(n3552), .Z(n3554) );
  HS65_LL_NOR2X3 U6537 ( .A(n4725), .B(n5422), .Z(n5499) );
  HS65_LH_AOI21X2 U6540 ( .A(n5192), .B(n5364), .C(n5500), .Z(n5365) );
  HS65_LH_IVX4 U6542 ( .A(n5271), .Z(n4246) );
  HS65_LL_NAND2X2 U6544 ( .A(n5516), .B(n5297), .Z(n5334) );
  HS65_LL_OAI12X3 U6545 ( .A(n5947), .B(n5950), .C(n5949), .Z(n6055) );
  HS65_LH_NAND2X4 U6546 ( .A(n4107), .B(n4106), .Z(n4111) );
  HS65_LH_IVX9 U6548 ( .A(n5342), .Z(n5569) );
  HS65_LH_NAND2X4 U6549 ( .A(\lte_x_59/B[21] ), .B(n4551), .Z(n3550) );
  HS65_LLS_XOR2X3 U6550 ( .A(n5951), .B(n2876), .Z(
        \u_DataPath/u_execute/resAdd1_i [29]) );
  HS65_LH_NAND2X4 U6552 ( .A(n4700), .B(n4699), .Z(n5356) );
  HS65_LH_OAI12X3 U6553 ( .A(n4425), .B(n4371), .C(n4373), .Z(n5606) );
  HS65_LH_NAND2X4 U6555 ( .A(n4701), .B(n5418), .Z(n5292) );
  HS65_LH_NOR2X3 U6559 ( .A(n5311), .B(n5299), .Z(n5540) );
  HS65_LH_NAND2X4 U6561 ( .A(\lte_x_59/B[5] ), .B(n4588), .Z(n3518) );
  HS65_LL_NOR2X3 U6562 ( .A(n4622), .B(n4630), .Z(n3491) );
  HS65_LH_NOR2X6 U6563 ( .A(n4880), .B(n4876), .Z(n4037) );
  HS65_LH_CNIVX3 U6564 ( .A(n5624), .Z(n3713) );
  HS65_LH_OAI12X3 U6566 ( .A(n5605), .B(n3731), .C(n3733), .Z(n3498) );
  HS65_LH_NAND2X4 U6569 ( .A(\lte_x_59/B[6] ), .B(n4544), .Z(n4462) );
  HS65_LH_OAI22X3 U6570 ( .A(n5179), .B(n2865), .C(n2848), .D(n4165), .Z(n4166) );
  HS65_LL_NOR2X2 U6571 ( .A(n5310), .B(n5095), .Z(n5552) );
  HS65_LH_IVX9 U6573 ( .A(n3575), .Z(n5192) );
  HS65_LH_OAI22X3 U6574 ( .A(n4682), .B(n4795), .C(n5129), .D(n5031), .Z(n4131) );
  HS65_LH_IVX9 U6575 ( .A(\sub_x_53/A[29] ), .Z(n4725) );
  HS65_LH_NAND2X4 U6576 ( .A(n4675), .B(n4674), .Z(n5517) );
  HS65_LH_NAND2X4 U6577 ( .A(n4663), .B(n3330), .Z(n4648) );
  HS65_LH_NAND2X4 U6578 ( .A(\lte_x_59/B[16] ), .B(n4587), .Z(n3910) );
  HS65_LH_NOR2X6 U6579 ( .A(\lte_x_59/B[15] ), .B(n5062), .Z(n3932) );
  HS65_LH_IVX9 U6580 ( .A(n4244), .Z(n5275) );
  HS65_LH_NAND2X7 U6581 ( .A(\lte_x_59/B[15] ), .B(n5062), .Z(n3934) );
  HS65_LH_NOR2X5 U6582 ( .A(n4341), .B(n4939), .Z(n4027) );
  HS65_LH_NOR2AX3 U6583 ( .A(n4587), .B(n2848), .Z(n3670) );
  HS65_LL_OAI12X2 U6586 ( .A(n4144), .B(n4481), .C(n4143), .Z(n4640) );
  HS65_LH_OAI12X3 U6587 ( .A(n4573), .B(n4570), .C(n4572), .Z(n3317) );
  HS65_LH_NAND2X4 U6588 ( .A(n4882), .B(n3855), .Z(n3856) );
  HS65_LH_CNIVX3 U6589 ( .A(n4081), .Z(n4082) );
  HS65_LH_NOR2X6 U6590 ( .A(n4371), .B(n4374), .Z(n5608) );
  HS65_LL_NOR2X3 U6592 ( .A(n3515), .B(n5530), .Z(n5271) );
  HS65_LH_IVX9 U6593 ( .A(n3814), .Z(n4051) );
  HS65_LH_CNIVX3 U6596 ( .A(n5503), .Z(n5504) );
  HS65_LL_NOR2X3 U6597 ( .A(n3846), .B(n4081), .Z(n4930) );
  HS65_LH_NAND2X2 U6599 ( .A(\lte_x_59/B[15] ), .B(n4588), .Z(n3644) );
  HS65_LL_AOI12X3 U6600 ( .A(\sub_x_53/A[27] ), .B(n3385), .C(n5343), .Z(n5582) );
  HS65_LH_IVX9 U6601 ( .A(n3560), .Z(n4845) );
  HS65_LH_NAND2X4 U6602 ( .A(\lte_x_59/B[14] ), .B(n4587), .Z(n4062) );
  HS65_LH_IVX9 U6604 ( .A(n5207), .Z(n5621) );
  HS65_LL_NOR2X2 U6606 ( .A(n3698), .B(n5627), .Z(n3379) );
  HS65_LH_OAI22X4 U6608 ( .A(n7917), .B(n8449), .C(n7916), .D(n8448), .Z(
        \u_DataPath/data_read_ex_1_i [29]) );
  HS65_LH_OAI22X4 U6609 ( .A(n7917), .B(n8415), .C(n7916), .D(n8414), .Z(
        \u_DataPath/data_read_ex_1_i [5]) );
  HS65_LH_OAI22X4 U6610 ( .A(n7917), .B(n8412), .C(n7916), .D(n8411), .Z(
        \u_DataPath/data_read_ex_1_i [20]) );
  HS65_LH_OAI22X4 U6611 ( .A(n7917), .B(n8457), .C(n7916), .D(n8455), .Z(
        \u_DataPath/data_read_ex_1_i [18]) );
  HS65_LH_OAI22X4 U6612 ( .A(n7917), .B(n8422), .C(n7916), .D(n8421), .Z(
        \u_DataPath/data_read_ex_1_i [31]) );
  HS65_LH_OAI22X4 U6613 ( .A(n7917), .B(n8408), .C(n7916), .D(n8407), .Z(
        \u_DataPath/data_read_ex_1_i [17]) );
  HS65_LH_OAI22X4 U6614 ( .A(n7917), .B(n7932), .C(n7916), .D(n8418), .Z(
        \u_DataPath/data_read_ex_1_i [28]) );
  HS65_LH_NOR2X6 U6615 ( .A(\lte_x_59/B[18] ), .B(n3371), .Z(n4244) );
  HS65_LH_NAND2X4 U6616 ( .A(n5130), .B(n5088), .Z(n5318) );
  HS65_LL_NAND2X4 U6617 ( .A(n5249), .B(n3788), .Z(n5624) );
  HS65_LL_NOR2AX3 U6621 ( .A(n2848), .B(n4147), .Z(n4630) );
  HS65_LH_NAND2X4 U6622 ( .A(n9188), .B(n9093), .Z(n7866) );
  HS65_LL_NAND2X4 U6627 ( .A(n4726), .B(n4966), .Z(n5572) );
  HS65_LH_NAND2X5 U6629 ( .A(n2849), .B(n5231), .Z(n5256) );
  HS65_LH_OAI21X3 U6630 ( .A(n3352), .B(n5179), .C(n4459), .Z(n4460) );
  HS65_LH_NAND2X4 U6631 ( .A(n2851), .B(n7627), .Z(n4229) );
  HS65_LH_NOR2X6 U6633 ( .A(\lte_x_59/B[21] ), .B(n3377), .Z(n4407) );
  HS65_LH_IVX9 U6634 ( .A(n3547), .Z(n4711) );
  HS65_LH_NAND2X4 U6635 ( .A(\sub_x_53/A[17] ), .B(n2870), .Z(n5531) );
  HS65_LL_AOI12X2 U6639 ( .A(n6117), .B(n6119), .C(n5943), .Z(n5950) );
  HS65_LL_NOR2X3 U6640 ( .A(\lte_x_59/B[5] ), .B(n4665), .Z(n4144) );
  HS65_LL_NOR2X5 U6641 ( .A(n4863), .B(n4838), .Z(n4887) );
  HS65_LH_NOR2X3 U6642 ( .A(n4147), .B(n2848), .Z(n5310) );
  HS65_LL_NOR2X3 U6643 ( .A(\lte_x_59/B[14] ), .B(n3366), .Z(n4913) );
  HS65_LH_NAND2X5 U6644 ( .A(\sub_x_53/A[23] ), .B(n5417), .Z(n5509) );
  HS65_LH_NOR4ABX2 U6645 ( .A(n6995), .B(n6994), .C(n6993), .D(n6992), .Z(
        n8338) );
  HS65_LH_NOR4ABX2 U6646 ( .A(n7035), .B(n7034), .C(n7033), .D(n7032), .Z(
        n8331) );
  HS65_LH_NOR4ABX2 U6647 ( .A(n7055), .B(n7054), .C(n7053), .D(n7052), .Z(
        n8327) );
  HS65_LH_NOR4ABX2 U6648 ( .A(n7075), .B(n7074), .C(n7073), .D(n7072), .Z(
        n8344) );
  HS65_LH_NOR4ABX2 U6649 ( .A(n7015), .B(n7014), .C(n7013), .D(n7012), .Z(
        n8349) );
  HS65_LH_NOR4ABX2 U6650 ( .A(n6361), .B(n6360), .C(n6359), .D(n6358), .Z(
        n8386) );
  HS65_LH_NOR4ABX2 U6651 ( .A(n6766), .B(n6765), .C(n6764), .D(n6763), .Z(
        n8322) );
  HS65_LL_NOR2X6 U6653 ( .A(n3151), .B(n3150), .Z(\lte_x_59/B[26] ) );
  HS65_LH_IVX9 U6655 ( .A(n5567), .Z(n3384) );
  HS65_LH_IVX9 U6656 ( .A(n5040), .Z(n4665) );
  HS65_LL_NAND2X4 U6660 ( .A(n8383), .B(n3237), .Z(n4969) );
  HS65_LHS_XOR2X3 U6665 ( .A(n5956), .B(n5955), .Z(
        \u_DataPath/u_execute/resAdd1_i [27]) );
  HS65_LL_OAI12X3 U6668 ( .A(n5748), .B(n5751), .C(n5750), .Z(n5908) );
  HS65_LH_OAI211X4 U6669 ( .A(n9243), .B(n8880), .C(n8295), .D(n9086), .Z(
        \u_DataPath/from_mem_data_out_i [10]) );
  HS65_LL_OAI12X2 U6672 ( .A(n8964), .B(n8088), .C(n8829), .Z(
        \u_DataPath/cw_to_ex_i [4]) );
  HS65_LL_OR2X9 U6674 ( .A(n3100), .B(n3099), .Z(n3101) );
  HS65_LH_NAND2X4 U6676 ( .A(n3352), .B(\lte_x_59/B[4] ), .Z(n5387) );
  HS65_LH_IVX9 U6677 ( .A(\sub_x_53/A[2] ), .Z(n5130) );
  HS65_LH_NAND2X7 U6678 ( .A(\lte_x_59/B[1] ), .B(n4805), .Z(n4824) );
  HS65_LH_NOR2X5 U6679 ( .A(\lte_x_59/B[3] ), .B(n5321), .Z(n3488) );
  HS65_LL_NOR2X6 U6680 ( .A(n3091), .B(n3090), .Z(\lte_x_59/B[14] ) );
  HS65_LH_NOR2X5 U6681 ( .A(n9167), .B(n8104), .Z(\u_DataPath/cw_to_ex_i [19])
         );
  HS65_LH_IVX7 U6682 ( .A(n5136), .Z(n5123) );
  HS65_LH_NAND2X4 U6683 ( .A(n5652), .B(n5654), .Z(n5362) );
  HS65_LL_IVX7 U6684 ( .A(\lte_x_59/B[8] ), .Z(n4682) );
  HS65_LL_OAI12X3 U6688 ( .A(n8176), .B(n3409), .C(n3408), .Z(n3410) );
  HS65_LH_AO22X9 U6689 ( .A(n8820), .B(n9138), .C(n9326), .D(n9153), .Z(
        \u_DataPath/jaddr_i [23]) );
  HS65_LL_NAND2X5 U6690 ( .A(n4191), .B(n4190), .Z(n7623) );
  HS65_LH_IVX9 U6691 ( .A(n5048), .Z(n3365) );
  HS65_LH_AO22X9 U6692 ( .A(n8819), .B(n9252), .C(n9327), .D(n9153), .Z(
        \u_DataPath/jaddr_i [24]) );
  HS65_LL_OAI22X3 U6693 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [19]), .C(
        n8323), .D(n3409), .Z(n3186) );
  HS65_LL_OAI22X3 U6695 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [18]), .C(
        n8387), .D(n3409), .Z(n3085) );
  HS65_LH_IVX4 U6696 ( .A(\u_DataPath/u_idexreg/N15 ), .Z(n8072) );
  HS65_LL_OAI12X6 U6697 ( .A(n3255), .B(n3254), .C(n3253), .Z(n4674) );
  HS65_LHS_XNOR2X3 U6698 ( .A(n7119), .B(n7122), .Z(
        \u_DataPath/u_execute/link_value_i [26]) );
  HS65_LL_OAI12X3 U6699 ( .A(n8389), .B(n3409), .C(n3089), .Z(n3090) );
  HS65_LL_NAND2AX7 U6700 ( .A(n2923), .B(n3281), .Z(n5061) );
  HS65_LH_AO22X9 U6702 ( .A(n8818), .B(n9252), .C(n9318), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [15]) );
  HS65_LH_IVX9 U6703 ( .A(n4534), .Z(n4431) );
  HS65_LL_NAND2AX7 U6709 ( .A(n3169), .B(n3168), .Z(n5652) );
  HS65_LH_AO22X9 U6711 ( .A(n8817), .B(n9138), .C(n9324), .D(n9153), .Z(
        \u_DataPath/jaddr_i [21]) );
  HS65_LH_AO22X9 U6712 ( .A(n8816), .B(n9138), .C(n9323), .D(n9153), .Z(
        \u_DataPath/jaddr_i [20]) );
  HS65_LL_NOR2X9 U6713 ( .A(n3316), .B(n3315), .Z(n5321) );
  HS65_LH_BFX18 U6715 ( .A(n9086), .Z(n7913) );
  HS65_LL_NAND2X5 U6716 ( .A(n3180), .B(n3179), .Z(n4699) );
  HS65_LH_OAI22X6 U6717 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [20]), .C(
        n8385), .D(n3409), .Z(n3176) );
  HS65_LH_AOI22X3 U6720 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ), .D(
        n7264), .Z(n6458) );
  HS65_LH_AO22X9 U6722 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ), .Z(n7361)
         );
  HS65_LH_AOI22X3 U6723 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][20] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ), .D(n7516), 
        .Z(n7479) );
  HS65_LH_AOI22X3 U6724 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ), .D(
        n2889), .Z(n7544) );
  HS65_LH_AOI22X3 U6726 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ), .D(n6942), .Z(n6487) );
  HS65_LH_AOI22X3 U6728 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ), .D(
        n2889), .Z(n7458) );
  HS65_LH_AOI22X3 U6730 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ), .D(
        n7264), .Z(n6478) );
  HS65_LH_AO22X9 U6731 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][6] ), .D(n7267), .Z(n6475) );
  HS65_LH_AOI22X3 U6733 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][8] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ), .D(n6942), .Z(n6467) );
  HS65_LH_AOI22X3 U6736 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ), .D(
        n2889), .Z(n7564) );
  HS65_LH_AOI22X3 U6737 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ), .D(
        n7264), .Z(n6558) );
  HS65_LH_AOI22X3 U6738 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ), .D(
        n2891), .Z(n7561) );
  HS65_LH_AOI22X3 U6739 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ), .D(n6942), .Z(n6567) );
  HS65_LH_AOI22X3 U6740 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][2] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ), .D(
        n6670), .Z(n6956) );
  HS65_LH_AOI22X3 U6742 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][19] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ), .D(
        n7264), .Z(n6518) );
  HS65_LH_AOI22X3 U6743 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ), .D(
        n6942), .Z(n6527) );
  HS65_LH_AO22X9 U6747 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][25] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ), .D(
        n7292), .Z(n7155) );
  HS65_LH_AOI22X3 U6748 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][25] ), .D(
        n6363), .Z(n7145) );
  HS65_LH_AOI22X3 U6750 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ), .D(n7516), 
        .Z(n6338) );
  HS65_LH_AO22X9 U6751 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ), .B(n7585), 
        .C(n6957), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ), .Z(n7411)
         );
  HS65_LH_AO22X9 U6752 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ), .D(n9372), .Z(n6597) );
  HS65_LH_AOI22X3 U6754 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ), .B(n7586), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][30] ), .D(
        n7587), .Z(n7414) );
  HS65_LH_AOI22X3 U6755 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ), .D(
        n7264), .Z(n6599) );
  HS65_LH_AOI22X3 U6756 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][10] ), .D(
        n7264), .Z(n6397) );
  HS65_LH_AOI22X3 U6758 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][7] ), .D(
        n7264), .Z(n6438) );
  HS65_LH_AOI22X3 U6759 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][7] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ), .D(n6942), .Z(n6447) );
  HS65_LH_AOI22X3 U6760 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ), .D(
        n7264), .Z(n6417) );
  HS65_LH_AOI22X3 U6761 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][12] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ), .D(
        n6942), .Z(n6547) );
  HS65_LH_AOI22X3 U6762 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ), .D(
        n7264), .Z(n6538) );
  HS65_LH_AOI22X3 U6764 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ), .D(n6942), .Z(n6609) );
  HS65_LH_AOI22X3 U6765 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ), .D(
        n6942), .Z(n6507) );
  HS65_LH_AOI22X3 U6766 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][0] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][0] ), .D(n6942), .Z(n6427) );
  HS65_LH_BFX18 U6767 ( .A(n8482), .Z(n7918) );
  HS65_LH_NAND2X7 U6771 ( .A(n8540), .B(n3178), .Z(n3179) );
  HS65_LL_NAND4ABX3 U6772 ( .A(n8558), .B(n4713), .C(n3146), .D(n8560), .Z(
        n3147) );
  HS65_LH_NOR2X5 U6773 ( .A(rst), .B(n8503), .Z(
        \u_DataPath/mem_writedata_out_i [8]) );
  HS65_LH_NAND2X5 U6776 ( .A(n7871), .B(n7870), .Z(
        \u_DataPath/mem_writedata_out_i [0]) );
  HS65_LH_AO22X9 U6780 ( .A(n9254), .B(n8815), .C(n9240), .D(n8984), .Z(
        \u_DataPath/pc4_to_idexreg_i [14]) );
  HS65_LH_AO22X9 U6781 ( .A(n9254), .B(n8814), .C(n9240), .D(n9097), .Z(
        \u_DataPath/pc4_to_idexreg_i [15]) );
  HS65_LH_AO22X9 U6782 ( .A(n9254), .B(n8813), .C(n9240), .D(n8979), .Z(
        \u_DataPath/pc4_to_idexreg_i [19]) );
  HS65_LH_IVX9 U6783 ( .A(n5032), .Z(n3352) );
  HS65_LH_AO22X9 U6784 ( .A(n9254), .B(n8812), .C(n9240), .D(n8985), .Z(
        \u_DataPath/pc4_to_idexreg_i [20]) );
  HS65_LL_IVX4 U6785 ( .A(n5030), .Z(n5312) );
  HS65_LL_OAI12X5 U6786 ( .A(n4216), .B(n4215), .C(n4214), .Z(n5422) );
  HS65_LH_NOR2X6 U6787 ( .A(n8846), .B(n3341), .Z(n3139) );
  HS65_LH_AO22X9 U6788 ( .A(n9254), .B(n8811), .C(n9273), .D(n9240), .Z(
        \u_DataPath/pc4_to_idexreg_i [2]) );
  HS65_LH_AO22X9 U6789 ( .A(n9254), .B(n8810), .C(n9240), .D(n8970), .Z(
        \u_DataPath/pc4_to_idexreg_i [3]) );
  HS65_LL_AOI12X4 U6790 ( .A(n3082), .B(n3335), .C(n3334), .Z(\lte_x_59/B[5] )
         );
  HS65_LH_AO22X9 U6791 ( .A(n9254), .B(n8809), .C(n9240), .D(n8971), .Z(
        \u_DataPath/pc4_to_idexreg_i [5]) );
  HS65_LH_AO22X9 U6792 ( .A(n9254), .B(n8808), .C(n8688), .D(n9240), .Z(
        \u_DataPath/pc4_to_idexreg_i [1]) );
  HS65_LH_AO22X9 U6794 ( .A(n9254), .B(n8806), .C(n9240), .D(n9098), .Z(
        \u_DataPath/pc4_to_idexreg_i [7]) );
  HS65_LH_AO22X9 U6795 ( .A(n9254), .B(n8805), .C(n9240), .D(n9010), .Z(
        \u_DataPath/pc4_to_idexreg_i [8]) );
  HS65_LL_OAI12X3 U6798 ( .A(n4210), .B(n2909), .C(n4209), .Z(n4966) );
  HS65_LH_AO22X9 U6802 ( .A(n9254), .B(n8803), .C(n9240), .D(n8981), .Z(
        \u_DataPath/pc4_to_idexreg_i [13]) );
  HS65_LH_IVX7 U6803 ( .A(n8053), .Z(n8054) );
  HS65_LH_IVX7 U6805 ( .A(n8059), .Z(\u_DataPath/cw_exmem_i [9]) );
  HS65_LH_NOR2AX6 U6806 ( .A(n3314), .B(n3414), .Z(n3316) );
  HS65_LH_NOR2X6 U6807 ( .A(n8858), .B(n3341), .Z(n3306) );
  HS65_LH_NOR2X6 U6808 ( .A(n8836), .B(n3341), .Z(n3061) );
  HS65_LL_NAND2X2 U6809 ( .A(n2927), .B(n8552), .Z(n3144) );
  HS65_LH_AO22X9 U6810 ( .A(n9254), .B(n8802), .C(n9240), .D(n8980), .Z(
        \u_DataPath/pc4_to_idexreg_i [25]) );
  HS65_LH_NAND2X7 U6811 ( .A(n3276), .B(n8523), .Z(n3277) );
  HS65_LH_NOR2X6 U6814 ( .A(n8856), .B(n3403), .Z(n3266) );
  HS65_LL_NAND3X2 U6815 ( .A(n3279), .B(n3280), .C(n8520), .Z(n3281) );
  HS65_LH_OR2X9 U6816 ( .A(\u_DataPath/data_read_ex_1_i [10]), .B(n3341), .Z(
        n3236) );
  HS65_LL_NOR2X3 U6817 ( .A(n3338), .B(n7863), .Z(n4657) );
  HS65_LH_NAND2AX7 U6818 ( .A(n8839), .B(n3291), .Z(n8548) );
  HS65_LH_NAND2AX7 U6820 ( .A(n8866), .B(n2874), .Z(n8545) );
  HS65_LL_NAND3X5 U6821 ( .A(n2879), .B(n8576), .C(n8318), .Z(n8401) );
  HS65_LL_NAND2X2 U6822 ( .A(n3221), .B(n5692), .Z(n3223) );
  HS65_LH_NAND2AX7 U6823 ( .A(\u_DataPath/data_read_ex_2_i [15]), .B(n2874), 
        .Z(n8523) );
  HS65_LL_NAND2AX4 U6824 ( .A(n3301), .B(n3300), .Z(n3302) );
  HS65_LH_NAND2AX7 U6825 ( .A(n8843), .B(n3291), .Z(n8532) );
  HS65_LL_NOR3X1 U6826 ( .A(n4713), .B(n8538), .C(n8539), .Z(n3178) );
  HS65_LH_NAND2AX7 U6827 ( .A(n8720), .B(n2874), .Z(n8540) );
  HS65_LL_NOR2X2 U6828 ( .A(n3154), .B(n8555), .Z(n3155) );
  HS65_LH_NAND2AX7 U6829 ( .A(n8721), .B(n3291), .Z(n8560) );
  HS65_LH_NAND2AX7 U6830 ( .A(n8832), .B(n2874), .Z(n8571) );
  HS65_LL_OAI22X3 U6832 ( .A(n3062), .B(n3340), .C(
        \u_DataPath/dataOut_exe_i [1]), .D(n3264), .Z(n3063) );
  HS65_LH_NAND2AX7 U6833 ( .A(n8718), .B(n3291), .Z(n8526) );
  HS65_LH_NAND2AX7 U6834 ( .A(n8837), .B(n3291), .Z(n8529) );
  HS65_LL_NAND2X7 U6835 ( .A(n2733), .B(n7902), .Z(n8443) );
  HS65_LL_AOI12X2 U6836 ( .A(n3142), .B(n2866), .C(n3141), .Z(n2927) );
  HS65_LL_NAND2X4 U6838 ( .A(n8703), .B(n7704), .Z(n7770) );
  HS65_LH_NAND2AX7 U6839 ( .A(n8717), .B(n2874), .Z(n8543) );
  HS65_LL_MUXI21X2 U6841 ( .D0(n8554), .D1(n4715), .S0(n4717), .Z(n3593) );
  HS65_LH_NAND2AX7 U6842 ( .A(n8865), .B(n2874), .Z(n8517) );
  HS65_LH_AOI22X4 U6843 ( .A(n8383), .B(n2866), .C(n3128), .D(n3291), .Z(n8561) );
  HS65_LH_NAND2AX7 U6844 ( .A(n8723), .B(n3291), .Z(n8520) );
  HS65_LH_NAND2X5 U6845 ( .A(n9084), .B(n8634), .Z(n8059) );
  HS65_LL_NOR2X5 U6846 ( .A(n3313), .B(n3312), .Z(n3414) );
  HS65_LL_NOR2X2 U6847 ( .A(n4188), .B(n8570), .Z(n4189) );
  HS65_LL_NOR2X2 U6848 ( .A(n3206), .B(n8525), .Z(n3207) );
  HS65_LH_NOR2X5 U6849 ( .A(n7673), .B(n7757), .Z(n7674) );
  HS65_LH_NOR2AX3 U6852 ( .A(n4714), .B(n5693), .Z(n3221) );
  HS65_LH_NAND2X7 U6853 ( .A(n3215), .B(n2896), .Z(n5691) );
  HS65_LH_NAND2X4 U6854 ( .A(n4714), .B(n8569), .Z(n2909) );
  HS65_LH_NOR2X5 U6855 ( .A(n3123), .B(n7671), .Z(n7672) );
  HS65_LH_NOR2X6 U6858 ( .A(n7657), .B(n7757), .Z(n7767) );
  HS65_LL_OAI12X12 U6859 ( .A(n3010), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N129 ) );
  HS65_LH_NAND2X4 U6861 ( .A(n4714), .B(n8565), .Z(n4215) );
  HS65_LL_OAI12X12 U6862 ( .A(n3009), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N92 ) );
  HS65_LH_NAND2X4 U6863 ( .A(n9376), .B(n8496), .Z(n3338) );
  HS65_LL_OAI12X12 U6864 ( .A(n8147), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N127 ) );
  HS65_LH_NOR2X6 U6865 ( .A(n7685), .B(n7757), .Z(n7764) );
  HS65_LH_NAND2X7 U6871 ( .A(n3278), .B(n3407), .Z(n3089) );
  HS65_LH_NAND2X4 U6872 ( .A(n4714), .B(n8533), .Z(n3194) );
  HS65_LL_NAND2X4 U6873 ( .A(n9376), .B(n8486), .Z(n3394) );
  HS65_LHS_XNOR2X6 U6874 ( .A(n5869), .B(n5868), .Z(\u_DataPath/toPC2_i [16])
         );
  HS65_LH_NAND2X4 U6875 ( .A(n7869), .B(n8621), .Z(n7871) );
  HS65_LH_NAND2X4 U6876 ( .A(n8235), .B(\u_DataPath/u_fetch/pc1/N3 ), .Z(n8044) );
  HS65_LL_NOR2X2 U6877 ( .A(n8488), .B(n9401), .Z(n3301) );
  HS65_LH_AND2X4 U6878 ( .A(\u_DataPath/dataOut_exe_i [15]), .B(n3407), .Z(
        n3271) );
  HS65_LH_NAND2X7 U6879 ( .A(n9376), .B(n8487), .Z(n3298) );
  HS65_LH_IVX7 U6880 ( .A(n8280), .Z(\u_DataPath/branch_target_i [4]) );
  HS65_LH_IVX7 U6881 ( .A(n8281), .Z(\u_DataPath/branch_target_i [3]) );
  HS65_LH_NAND2X4 U6882 ( .A(n9376), .B(n8502), .Z(n3329) );
  HS65_LHS_XNOR2X6 U6883 ( .A(n7732), .B(n7731), .Z(
        \u_DataPath/u_execute/link_value_i [13]) );
  HS65_LHS_XNOR2X6 U6884 ( .A(n7722), .B(n7721), .Z(
        \u_DataPath/u_execute/link_value_i [15]) );
  HS65_LH_IVX18 U6885 ( .A(n4548), .Z(n5648) );
  HS65_LH_AOI12X2 U6887 ( .A(n6069), .B(n6071), .C(n5984), .Z(n5985) );
  HS65_LHS_XNOR2X6 U6888 ( .A(n6080), .B(n6079), .Z(
        \u_DataPath/u_execute/resAdd1_i [9]) );
  HS65_LL_NAND2AX4 U6889 ( .A(n3034), .B(n3033), .Z(n3045) );
  HS65_LL_NAND2X7 U6890 ( .A(n2733), .B(n8160), .Z(n8117) );
  HS65_LH_AOI12X2 U6891 ( .A(n6002), .B(n6083), .C(n6001), .Z(n6003) );
  HS65_LHS_XNOR2X6 U6893 ( .A(n6084), .B(n6083), .Z(
        \u_DataPath/u_execute/resAdd1_i [16]) );
  HS65_LH_OAI12X3 U6894 ( .A(n5983), .B(n6077), .C(n5982), .Z(n6071) );
  HS65_LH_NOR2X5 U6895 ( .A(n5700), .B(n7710), .Z(n5701) );
  HS65_LH_IVX9 U6896 ( .A(n7653), .Z(n7749) );
  HS65_LH_NOR2X5 U6897 ( .A(n7711), .B(n7710), .Z(n7712) );
  HS65_LH_NAND2X5 U6898 ( .A(n3160), .B(n7802), .Z(n8549) );
  HS65_LH_OAI12X3 U6899 ( .A(n5964), .B(n6077), .C(n5963), .Z(n5992) );
  HS65_LH_NOR2X3 U6900 ( .A(n8847), .B(n7802), .Z(n3337) );
  HS65_LL_NAND2X5 U6901 ( .A(n3131), .B(n3217), .Z(n3310) );
  HS65_LL_NOR2AX3 U6902 ( .A(n3032), .B(n8262), .Z(n3033) );
  HS65_LH_OAI12X3 U6903 ( .A(n6078), .B(n6077), .C(n6076), .Z(n6079) );
  HS65_LH_OAI12X3 U6904 ( .A(n5782), .B(n5878), .C(n5781), .Z(n5872) );
  HS65_LL_NAND2X5 U6905 ( .A(n3217), .B(n3131), .Z(n2896) );
  HS65_LH_OAI12X3 U6906 ( .A(n5879), .B(n5878), .C(n5877), .Z(n5880) );
  HS65_LH_NOR2X3 U6909 ( .A(n8092), .B(n7762), .Z(n8075) );
  HS65_LL_OAI12X3 U6910 ( .A(n5939), .B(n5999), .C(n5938), .Z(n6111) );
  HS65_LH_NAND2X4 U6911 ( .A(n9114), .B(n9369), .Z(n8429) );
  HS65_LH_IVX4 U6912 ( .A(n7692), .Z(n7682) );
  HS65_LHS_XNOR2X6 U6913 ( .A(n5893), .B(n5892), .Z(\u_DataPath/toPC2_i [4])
         );
  HS65_LL_NOR4ABX9 U6914 ( .A(n2954), .B(n2953), .C(n2952), .D(n2951), .Z(
        n3217) );
  HS65_LL_NAND2X4 U6915 ( .A(n3057), .B(n3028), .Z(n2932) );
  HS65_LH_NOR2X6 U6917 ( .A(n7834), .B(n3442), .Z(n3431) );
  HS65_LHS_XNOR2X6 U6918 ( .A(n2835), .B(n7746), .Z(\u_DataPath/pc_4_i [8]) );
  HS65_LH_IVX7 U6919 ( .A(n7684), .Z(n7685) );
  HS65_LH_AOI21X6 U6920 ( .A(n5934), .B(n5962), .C(n5933), .Z(n5999) );
  HS65_LH_NAND3X5 U6921 ( .A(n7698), .B(n7697), .C(n7777), .Z(n8083) );
  HS65_LL_AOI12X2 U6922 ( .A(n6013), .B(n6015), .C(n5937), .Z(n5938) );
  HS65_LH_NAND2X5 U6924 ( .A(n7091), .B(n7090), .Z(n7092) );
  HS65_LL_NAND2X2 U6925 ( .A(n9111), .B(n3049), .Z(n3051) );
  HS65_LH_NOR2X3 U6926 ( .A(n8086), .B(n8098), .Z(n7762) );
  HS65_LH_NOR2X5 U6929 ( .A(n7788), .B(n7787), .Z(n7708) );
  HS65_LH_NAND2X4 U6930 ( .A(n3395), .B(n5716), .Z(n3398) );
  HS65_LL_NOR2X2 U6932 ( .A(n3048), .B(n3054), .Z(n3032) );
  HS65_LH_NAND3X3 U6933 ( .A(n3011), .B(n9076), .C(n9078), .Z(n3012) );
  HS65_LH_OAI12X3 U6934 ( .A(n5899), .B(n5898), .C(n5897), .Z(n5900) );
  HS65_LHS_XOR2X6 U6935 ( .A(n8943), .B(n2846), .Z(n3028) );
  HS65_LL_NAND2X4 U6936 ( .A(n2945), .B(n2944), .Z(n2954) );
  HS65_LL_NOR2AX3 U6937 ( .A(n2733), .B(n5716), .Z(n7861) );
  HS65_LL_NOR2X5 U6938 ( .A(n6348), .B(n6341), .Z(n6680) );
  HS65_LH_NOR2X5 U6939 ( .A(n8090), .B(n7700), .Z(n8097) );
  HS65_LL_NOR2X5 U6940 ( .A(n6148), .B(n6140), .Z(n6171) );
  HS65_LL_NOR2X5 U6941 ( .A(n6350), .B(n6341), .Z(n6754) );
  HS65_LH_NOR2X5 U6942 ( .A(n7742), .B(n7741), .Z(n7666) );
  HS65_LH_OAI12X3 U6944 ( .A(n6102), .B(n6101), .C(n6100), .Z(n6103) );
  HS65_LL_NOR2X5 U6945 ( .A(n6146), .B(n6140), .Z(n6172) );
  HS65_LH_NAND2X4 U6946 ( .A(n5769), .B(n5768), .Z(n5771) );
  HS65_LH_NOR3X4 U6947 ( .A(n9233), .B(n8236), .C(rst), .Z(n8285) );
  HS65_LL_AOI21X2 U6948 ( .A(n5981), .B(n5928), .C(n5927), .Z(n5963) );
  HS65_LH_NAND2X4 U6949 ( .A(n5826), .B(n5825), .Z(n5828) );
  HS65_LH_NAND2X4 U6950 ( .A(n5750), .B(n5749), .Z(n5752) );
  HS65_LH_NAND2X4 U6951 ( .A(n6082), .B(n6081), .Z(n6084) );
  HS65_LH_NOR3X4 U6952 ( .A(n9236), .B(n9237), .C(n7638), .Z(n8269) );
  HS65_LH_NAND2X4 U6953 ( .A(n5788), .B(n5787), .Z(n5794) );
  HS65_LH_NOR2X5 U6954 ( .A(n2975), .B(n7638), .Z(n2978) );
  HS65_LH_IVX7 U6955 ( .A(n8115), .Z(n8123) );
  HS65_LL_NOR2X3 U6959 ( .A(n6349), .B(n2878), .Z(n6670) );
  HS65_LL_NOR2X5 U6960 ( .A(n6150), .B(n6151), .Z(n2888) );
  HS65_LH_NAND2X4 U6961 ( .A(n6075), .B(n5875), .Z(n6080) );
  HS65_LH_NAND2X4 U6962 ( .A(n5973), .B(n5972), .Z(n5975) );
  HS65_LL_NOR2X3 U6965 ( .A(n6350), .B(n6332), .Z(n6740) );
  HS65_LH_NAND2X4 U6966 ( .A(n6028), .B(n6027), .Z(n6030) );
  HS65_LH_NAND2X4 U6968 ( .A(n6100), .B(n6050), .Z(n6052) );
  HS65_LH_NAND2X4 U6969 ( .A(n4717), .B(n9343), .Z(n4214) );
  HS65_LH_NAND2X4 U6970 ( .A(n5954), .B(n5953), .Z(n5956) );
  HS65_LH_NAND2X4 U6972 ( .A(n4717), .B(n9341), .Z(n4970) );
  HS65_LL_NOR2X5 U6973 ( .A(n6348), .B(n6332), .Z(n6747) );
  HS65_LH_NAND3X5 U6974 ( .A(n2847), .B(n3008), .C(n7086), .Z(n3009) );
  HS65_LH_IVX7 U6976 ( .A(n5965), .Z(n5966) );
  HS65_LHS_XNOR2X6 U6977 ( .A(n7669), .B(n7743), .Z(\u_DataPath/pc_4_i [4]) );
  HS65_LHS_XNOR2X3 U6978 ( .A(n7726), .B(n7789), .Z(
        \u_DataPath/u_execute/link_value_i [4]) );
  HS65_LH_NAND2X4 U6979 ( .A(n4713), .B(n9341), .Z(n3204) );
  HS65_LH_NAND2X4 U6980 ( .A(n6094), .B(n5890), .Z(n6096) );
  HS65_LL_NOR2X5 U6981 ( .A(n6148), .B(n6139), .Z(n2887) );
  HS65_LL_NAND2AX4 U6983 ( .A(n3039), .B(n3038), .Z(n3042) );
  HS65_LH_MUXI21X2 U6985 ( .D0(n3406), .D1(n9395), .S0(n3404), .Z(n8176) );
  HS65_LH_NAND3X5 U6986 ( .A(n9237), .B(n2975), .C(n2973), .Z(n2974) );
  HS65_LH_NOR2X6 U6987 ( .A(n3121), .B(n7686), .Z(n7659) );
  HS65_LL_NAND2X4 U6989 ( .A(\u_DataPath/jaddr_i [24]), .B(n6126), .Z(n6151)
         );
  HS65_LH_NOR2X6 U6990 ( .A(\u_DataPath/jaddr_i [24]), .B(n8165), .Z(n6138) );
  HS65_LL_OR3X4 U6991 ( .A(n8165), .B(n8151), .C(\u_DataPath/jaddr_i [25]), 
        .Z(n6147) );
  HS65_LH_NOR2X5 U6992 ( .A(n8162), .B(n8074), .Z(n8086) );
  HS65_LLS_XNOR2X3 U6993 ( .A(n8944), .B(n8170), .Z(n3040) );
  HS65_LL_NAND2X4 U6994 ( .A(\u_DataPath/jaddr_i [25]), .B(n6145), .Z(n6139)
         );
  HS65_LH_NAND2X4 U6995 ( .A(n6118), .B(n6117), .Z(n6120) );
  HS65_LHS_XNOR2X3 U6996 ( .A(n9116), .B(n7706), .Z(
        \u_DataPath/u_execute/link_value_i [3]) );
  HS65_LH_MUXI21X2 U6997 ( .D0(n2956), .D1(n9394), .S0(n3404), .Z(n8364) );
  HS65_LH_NOR2X3 U6998 ( .A(\u_DataPath/immediate_ext_dec_i [3]), .B(n8090), 
        .Z(n8121) );
  HS65_LH_IVX4 U6999 ( .A(n8159), .Z(n8625) );
  HS65_LH_NAND3X5 U7000 ( .A(n9082), .B(n9068), .C(n7642), .Z(n7688) );
  HS65_LH_NAND2X5 U7001 ( .A(opcode_i[5]), .B(n7695), .Z(n8037) );
  HS65_LH_NOR2X3 U7004 ( .A(n8151), .B(rst), .Z(\u_DataPath/rs_ex_i [3]) );
  HS65_LH_NAND3X3 U7005 ( .A(n9082), .B(n7696), .C(n7695), .Z(n8041) );
  HS65_LH_NOR2X5 U7007 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .B(n8162), 
        .Z(n8096) );
  HS65_LL_MUXI21X2 U7008 ( .D0(n3212), .D1(n9396), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8265) );
  HS65_LH_NAND2X4 U7009 ( .A(n6114), .B(n6113), .Z(n6116) );
  HS65_LH_IVX4 U7011 ( .A(n5855), .Z(n5718) );
  HS65_LH_NAND2X4 U7013 ( .A(n5915), .B(n5914), .Z(n5917) );
  HS65_LH_NAND2X4 U7016 ( .A(n5911), .B(n5910), .Z(n5913) );
  HS65_LH_NOR2X6 U7017 ( .A(n7834), .B(n5491), .Z(n3421) );
  HS65_LH_OAI12X3 U7018 ( .A(n6006), .B(n5987), .C(n5989), .Z(n5965) );
  HS65_LL_NAND2X5 U7019 ( .A(n3030), .B(n2946), .Z(n3008) );
  HS65_LL_NAND3X2 U7020 ( .A(\u_DataPath/cw_to_ex_i [4]), .B(n5492), .C(n5491), 
        .Z(n5493) );
  HS65_LH_OAI12X3 U7021 ( .A(n6064), .B(n2875), .C(n6063), .Z(n5935) );
  HS65_LH_NOR2X5 U7023 ( .A(n5836), .B(n5839), .Z(n5834) );
  HS65_LH_NOR2X6 U7024 ( .A(n6085), .B(n6090), .Z(n5924) );
  HS65_LL_OAI12X2 U7025 ( .A(n5850), .B(n5846), .C(n5848), .Z(n5844) );
  HS65_LH_OAI12X3 U7026 ( .A(n6088), .B(n6085), .C(n6087), .Z(n5923) );
  HS65_LH_NAND2X4 U7027 ( .A(n5907), .B(n5906), .Z(n5909) );
  HS65_LL_NAND2AX7 U7029 ( .A(n9078), .B(n3030), .Z(n7084) );
  HS65_LH_OAI12X3 U7030 ( .A(n6076), .B(n6073), .C(n6075), .Z(n5981) );
  HS65_LH_IVX7 U7031 ( .A(n5867), .Z(n5821) );
  HS65_LH_NAND2AX7 U7032 ( .A(n8480), .B(n9347), .Z(n8051) );
  HS65_LH_NOR2X5 U7033 ( .A(n8942), .B(n9222), .Z(n6022) );
  HS65_LH_NOR2X3 U7034 ( .A(\u_DataPath/jaddr_i [23]), .B(
        \u_DataPath/jaddr_i [25]), .Z(n6126) );
  HS65_LH_MUX21X4 U7035 ( .D0(n8908), .D1(\u_DataPath/from_mem_data_out_i [6]), 
        .S0(\u_DataPath/cw_towb_i [0]), .Z(n8311) );
  HS65_LH_NOR2X3 U7036 ( .A(opcode_i[5]), .B(n9068), .Z(n7735) );
  HS65_LH_NOR2X5 U7039 ( .A(\u_DataPath/jaddr_i [18]), .B(
        \u_DataPath/jaddr_i [19]), .Z(n6339) );
  HS65_LH_NOR2X5 U7040 ( .A(n9342), .B(n9209), .Z(n5767) );
  HS65_LH_NOR2X5 U7041 ( .A(n9341), .B(n9213), .Z(n5824) );
  HS65_LH_NOR2X3 U7042 ( .A(\u_DataPath/immediate_ext_dec_i [5]), .B(
        \u_DataPath/immediate_ext_dec_i [4]), .Z(n8120) );
  HS65_LL_NOR2X3 U7043 ( .A(n9341), .B(n9221), .Z(n5817) );
  HS65_LH_NOR2X5 U7044 ( .A(n9341), .B(n9222), .Z(n5820) );
  HS65_LH_IVX9 U7046 ( .A(n7835), .Z(n7116) );
  HS65_LH_NAND2X4 U7047 ( .A(\u_DataPath/immediate_ext_dec_i [5]), .B(
        \u_DataPath/immediate_ext_dec_i [4]), .Z(n8074) );
  HS65_LH_NOR2X5 U7053 ( .A(n9175), .B(n9227), .Z(n5882) );
  HS65_LH_NOR2X3 U7054 ( .A(n9037), .B(n9212), .Z(n6045) );
  HS65_LLS_XNOR2X3 U7055 ( .A(n8761), .B(n9004), .Z(n3036) );
  HS65_LH_NAND2X7 U7056 ( .A(n9179), .B(n9225), .Z(n6088) );
  HS65_LH_NAND2X7 U7057 ( .A(n9175), .B(n9227), .Z(n6087) );
  HS65_LLS_XNOR2X3 U7058 ( .A(n8763), .B(n8942), .Z(n2960) );
  HS65_LLS_XNOR2X3 U7059 ( .A(n9077), .B(n8761), .Z(n2957) );
  HS65_LLS_XNOR2X3 U7060 ( .A(n8764), .B(n8967), .Z(n2963) );
  HS65_LH_IVX9 U7061 ( .A(n8762), .Z(n8107) );
  HS65_LH_NAND2X7 U7062 ( .A(n9177), .B(n9229), .Z(n6076) );
  HS65_LH_NAND2X7 U7064 ( .A(n9171), .B(n9214), .Z(n6070) );
  HS65_LL_OAI21X2 U7065 ( .A(\u_DataPath/cw_towb_i [1]), .B(n9075), .C(n9077), 
        .Z(n2944) );
  HS65_LL_IVX7 U7066 ( .A(n9076), .Z(n2946) );
  HS65_LH_NAND2X7 U7067 ( .A(n9232), .B(n9214), .Z(n7728) );
  HS65_LH_NAND2X7 U7068 ( .A(n9267), .B(n9228), .Z(n5989) );
  HS65_LH_NAND2X4 U7070 ( .A(n9342), .B(n9202), .Z(n5852) );
  HS65_LH_NOR2X5 U7071 ( .A(n9343), .B(n9203), .Z(n5855) );
  HS65_LH_NOR2X5 U7072 ( .A(n9145), .B(n9224), .Z(n5957) );
  HS65_LH_NOR2X5 U7073 ( .A(n9343), .B(n9205), .Z(n5743) );
  HS65_LH_NOR2X5 U7074 ( .A(n8968), .B(n9217), .Z(n5995) );
  HS65_LH_NOR2X6 U7075 ( .A(n8966), .B(n9221), .Z(n6019) );
  HS65_LH_OR2X9 U7076 ( .A(n9342), .B(n9206), .Z(n5906) );
  HS65_LH_NAND2X7 U7077 ( .A(n8966), .B(n9221), .Z(n6021) );
  HS65_LH_NOR2X5 U7078 ( .A(n9179), .B(n9225), .Z(n5887) );
  HS65_LH_NAND3X5 U7079 ( .A(opcode_i[3]), .B(opcode_i[5]), .C(n9068), .Z(
        n7636) );
  HS65_LH_IVX9 U7080 ( .A(n9113), .Z(n2983) );
  HS65_LL_NOR2X3 U7081 ( .A(n9237), .B(n8915), .Z(n2976) );
  HS65_LL_NAND3AX6 U7083 ( .A(n4833), .B(n4832), .C(n7848), .Z(n5679) );
  HS65_LL_NAND3AX3 U7084 ( .A(n5602), .B(n8479), .C(n8458), .Z(n5676) );
  HS65_LL_IVX4 U7086 ( .A(n5710), .Z(n5711) );
  HS65_LL_NOR2AX3 U7087 ( .A(n5709), .B(n5708), .Z(n7859) );
  HS65_LH_OAI12X3 U7088 ( .A(n9190), .B(n8888), .C(n8294), .Z(
        \u_DataPath/dataOut_exe_i [10]) );
  HS65_LH_NAND2X4 U7089 ( .A(n5285), .B(n5707), .Z(n4370) );
  HS65_LL_AO12X4 U7091 ( .A(n5285), .B(n5222), .C(n5221), .Z(n5224) );
  HS65_LL_NAND2AX4 U7092 ( .A(n4961), .B(n4960), .Z(n4962) );
  HS65_LH_NAND3X3 U7093 ( .A(n5704), .B(n8462), .C(n4537), .Z(n4833) );
  HS65_LL_NAND2AX4 U7094 ( .A(n3626), .B(n3625), .Z(n3627) );
  HS65_LH_CBI4I1X5 U7095 ( .A(n8883), .B(n9201), .C(n9239), .D(n7836), .Z(
        \u_DataPath/dataOut_exe_i [11]) );
  HS65_LH_AND2X9 U7096 ( .A(n5285), .B(n7626), .Z(n5598) );
  HS65_LHS_XNOR2X6 U7099 ( .A(n2915), .B(n4313), .Z(n5707) );
  HS65_LLS_XNOR2X3 U7101 ( .A(n2914), .B(n4300), .Z(n4301) );
  HS65_LL_AO12X4 U7102 ( .A(n4367), .B(n5285), .C(n4366), .Z(n4368) );
  HS65_LLS_XNOR2X3 U7103 ( .A(n4413), .B(n4412), .Z(n4414) );
  HS65_LLS_XNOR2X3 U7105 ( .A(n3580), .B(n3579), .Z(n3628) );
  HS65_LL_AO12X4 U7106 ( .A(n5643), .B(n4450), .C(n4449), .Z(n4451) );
  HS65_LHS_XNOR2X6 U7107 ( .A(n4935), .B(n4934), .Z(n4936) );
  HS65_LL_NOR3X1 U7108 ( .A(n5705), .B(n4536), .C(n6121), .Z(n4537) );
  HS65_LH_NOR2AX3 U7110 ( .A(n3799), .B(n3798), .Z(n3811) );
  HS65_LL_AND3X4 U7111 ( .A(n4901), .B(n4900), .C(n4899), .Z(n4910) );
  HS65_LL_NAND2X2 U7113 ( .A(n5217), .B(n4327), .Z(n4369) );
  HS65_LH_NAND2X7 U7115 ( .A(n5643), .B(n3566), .Z(n3567) );
  HS65_LLS_XNOR2X3 U7116 ( .A(n4242), .B(n4241), .Z(n7626) );
  HS65_LL_NAND2X2 U7117 ( .A(n4448), .B(n4447), .Z(n4449) );
  HS65_LL_AND3X4 U7118 ( .A(n5368), .B(n5341), .C(n5340), .Z(n2920) );
  HS65_LH_NAND2AX7 U7119 ( .A(n3797), .B(n3796), .Z(n3798) );
  HS65_LL_OAI21X3 U7120 ( .A(n4246), .B(n5633), .C(n4245), .Z(n4247) );
  HS65_LLS_XNOR2X3 U7122 ( .A(n4379), .B(n4378), .Z(n4380) );
  HS65_LLS_XNOR2X3 U7123 ( .A(n2907), .B(n9338), .Z(n3902) );
  HS65_LL_NAND2AX4 U7124 ( .A(n5076), .B(n5075), .Z(n5077) );
  HS65_LL_OAI12X3 U7125 ( .A(n5277), .B(n5633), .C(n5276), .Z(n5278) );
  HS65_LHS_XNOR2X6 U7126 ( .A(n3623), .B(n3622), .Z(n3624) );
  HS65_LL_OAI12X3 U7127 ( .A(n5633), .B(n4337), .C(n4336), .Z(n4338) );
  HS65_LL_NOR2AX3 U7128 ( .A(n4933), .B(n4932), .Z(n4934) );
  HS65_LLS_XNOR2X3 U7129 ( .A(n4226), .B(n4225), .Z(n7622) );
  HS65_LH_CBI4I1X5 U7130 ( .A(n8882), .B(n8894), .C(n9189), .D(n8436), .Z(
        \u_DataPath/dataOut_exe_i [2]) );
  HS65_LH_OAI21X3 U7131 ( .A(n3578), .B(n5633), .C(n3577), .Z(n3579) );
  HS65_LL_OAI12X3 U7132 ( .A(n4311), .B(n5633), .C(n4310), .Z(n4312) );
  HS65_LH_NAND2AX7 U7133 ( .A(n5593), .B(n5592), .Z(n5594) );
  HS65_LL_OAI12X3 U7134 ( .A(n4411), .B(n5633), .C(n4410), .Z(n4412) );
  HS65_LL_OAI12X3 U7135 ( .A(n5197), .B(n5633), .C(n5196), .Z(n5198) );
  HS65_LL_NAND3AX3 U7136 ( .A(n4172), .B(n4171), .C(n4170), .Z(n4173) );
  HS65_LL_NAND2X2 U7137 ( .A(n5339), .B(n5338), .Z(n5340) );
  HS65_LL_OAI12X3 U7138 ( .A(n5213), .B(n2859), .C(n5212), .Z(n5214) );
  HS65_LL_NAND2X2 U7139 ( .A(n5372), .B(n5371), .Z(n5596) );
  HS65_LL_NAND2AX4 U7140 ( .A(n3467), .B(n3466), .Z(n3468) );
  HS65_LHS_XNOR2X6 U7142 ( .A(n3943), .B(n3942), .Z(n3944) );
  HS65_LHS_XNOR2X6 U7143 ( .A(n3994), .B(n3993), .Z(n3995) );
  HS65_LL_AO12X4 U7144 ( .A(n5074), .B(n5073), .C(n5072), .Z(n5075) );
  HS65_LL_OAI12X3 U7145 ( .A(n3473), .B(n2859), .C(n4251), .Z(n4252) );
  HS65_LL_OAI12X3 U7146 ( .A(n5263), .B(n2859), .C(n5262), .Z(n5264) );
  HS65_LL_NOR2AX3 U7147 ( .A(n5591), .B(n5590), .Z(n5592) );
  HS65_LL_NAND3X2 U7148 ( .A(n4278), .B(n4277), .C(n4276), .Z(n4279) );
  HS65_LLS_XNOR2X3 U7149 ( .A(n4923), .B(n4922), .Z(n4963) );
  HS65_LL_NAND2AX4 U7151 ( .A(n5669), .B(n5668), .Z(n5670) );
  HS65_LL_NAND3AX3 U7152 ( .A(n3730), .B(n3729), .C(n3728), .Z(n3744) );
  HS65_LLS_XNOR2X3 U7153 ( .A(n2906), .B(n3817), .Z(n3852) );
  HS65_LL_OAI21X2 U7155 ( .A(n5152), .B(n4473), .C(n4472), .Z(n4474) );
  HS65_LL_NOR2AX3 U7156 ( .A(n4388), .B(n5152), .Z(n4122) );
  HS65_LL_NAND4X4 U7158 ( .A(n4567), .B(n4566), .C(n4565), .D(n4564), .Z(n4568) );
  HS65_LL_AOI21X2 U7159 ( .A(n3751), .B(n5195), .C(n3750), .Z(n3752) );
  HS65_LL_NAND2AX4 U7162 ( .A(n4520), .B(n4519), .Z(n4948) );
  HS65_LL_NAND2X2 U7163 ( .A(n5589), .B(n5588), .Z(n5590) );
  HS65_LL_OR3X4 U7164 ( .A(n4860), .B(n4859), .C(n4858), .Z(n2902) );
  HS65_LL_NAND3AX3 U7165 ( .A(n3929), .B(n3928), .C(n3927), .Z(n3930) );
  HS65_LH_OAI12X3 U7166 ( .A(n4387), .B(n4386), .C(n5672), .Z(n4406) );
  HS65_LL_NAND3X2 U7167 ( .A(n5112), .B(n5111), .C(n5110), .Z(n5113) );
  HS65_LL_NAND3X2 U7168 ( .A(n4152), .B(n4151), .C(n4150), .Z(n4172) );
  HS65_LL_NAND3AX3 U7169 ( .A(n3787), .B(n3786), .C(n3785), .Z(n3794) );
  HS65_LH_AOI21X2 U7170 ( .A(n5624), .B(n5623), .C(n5622), .Z(n5625) );
  HS65_LL_AOI22X1 U7171 ( .A(n6123), .B(n5250), .C(n4512), .D(n5248), .Z(n8462) );
  HS65_LL_AOI21X2 U7174 ( .A(n4222), .B(n5211), .C(n4221), .Z(n4223) );
  HS65_LL_NAND3X2 U7175 ( .A(n5584), .B(n5536), .C(n5535), .Z(n5537) );
  HS65_LH_OA12X4 U7176 ( .A(n3894), .B(n3815), .C(n3816), .Z(n3817) );
  HS65_LH_NOR4ABX2 U7177 ( .A(n5335), .B(n4017), .C(n5334), .D(n5333), .Z(
        n5336) );
  HS65_LH_OAI21X3 U7178 ( .A(n3981), .B(n5152), .C(n3980), .Z(n3988) );
  HS65_LH_NAND3X3 U7179 ( .A(n3655), .B(n3429), .C(n3428), .Z(n3467) );
  HS65_LL_NAND3X2 U7181 ( .A(n4980), .B(n4979), .C(n4978), .Z(n4995) );
  HS65_LL_CB4I1X4 U7182 ( .A(n4695), .B(n4694), .C(n4693), .D(n4692), .Z(n4784) );
  HS65_LH_OAI21X3 U7184 ( .A(n5646), .B(n4849), .C(n4848), .Z(n4860) );
  HS65_LH_AOI21X2 U7185 ( .A(n5207), .B(n5206), .C(n5205), .Z(n5219) );
  HS65_LH_AOI21X2 U7186 ( .A(n5659), .B(n5239), .C(n3675), .Z(n3676) );
  HS65_LL_NAND4ABX3 U7187 ( .A(n4621), .B(n4620), .C(n4619), .D(n4618), .Z(
        n4652) );
  HS65_LH_NAND3X3 U7188 ( .A(n3655), .B(n3654), .C(n3653), .Z(n3680) );
  HS65_LH_OAI21X3 U7189 ( .A(n4753), .B(n5656), .C(n4135), .Z(n4136) );
  HS65_LH_NAND3X3 U7190 ( .A(n4431), .B(n5089), .C(n4430), .Z(n4448) );
  HS65_LH_OAI21X3 U7191 ( .A(n4812), .B(n4811), .C(n4810), .Z(n4813) );
  HS65_LL_NAND2X2 U7192 ( .A(n4518), .B(n4517), .Z(n4520) );
  HS65_LH_OAI21X3 U7193 ( .A(n5177), .B(n5176), .C(n5175), .Z(n5190) );
  HS65_LH_NAND2X4 U7195 ( .A(n4309), .B(n5194), .Z(n4311) );
  HS65_LL_AOI12X2 U7196 ( .A(n4516), .B(n4515), .C(n4514), .Z(n4518) );
  HS65_LLS_XOR2X3 U7198 ( .A(n4104), .B(n4103), .Z(n4141) );
  HS65_LL_NAND3X2 U7199 ( .A(n4202), .B(n4201), .C(n4200), .Z(n4203) );
  HS65_LL_NAND2X2 U7200 ( .A(n5352), .B(n5351), .Z(n5482) );
  HS65_LL_OR2X4 U7201 ( .A(n3894), .B(n3370), .Z(n2929) );
  HS65_LH_NOR2AX3 U7203 ( .A(n5058), .B(n5057), .Z(n5059) );
  HS65_LL_NAND3X2 U7204 ( .A(n5297), .B(n5109), .C(n5108), .Z(n5526) );
  HS65_LLS_XOR2X3 U7205 ( .A(n4146), .B(n4145), .Z(n4174) );
  HS65_LH_IVX9 U7206 ( .A(n4918), .Z(n3816) );
  HS65_LH_AOI21X2 U7207 ( .A(n4951), .B(n4875), .C(n4874), .Z(n4901) );
  HS65_LH_NAND2X4 U7209 ( .A(n4007), .B(n4836), .Z(n4606) );
  HS65_LLS_XOR2X3 U7211 ( .A(n4648), .B(n4647), .Z(n4649) );
  HS65_LH_AOI21X2 U7212 ( .A(n3778), .B(n5658), .C(n3777), .Z(n3786) );
  HS65_LH_AOI21X2 U7213 ( .A(n5234), .B(n4033), .C(n4032), .Z(n4048) );
  HS65_LH_AOI21X2 U7214 ( .A(n5131), .B(n4615), .C(n4026), .Z(n2931) );
  HS65_LL_NOR2AX6 U7215 ( .A(n3482), .B(n3481), .Z(n3618) );
  HS65_LH_AOI21X2 U7216 ( .A(n5144), .B(n4560), .C(n4559), .Z(n4565) );
  HS65_LH_CNIVX3 U7219 ( .A(n5174), .Z(n3462) );
  HS65_LH_AOI21X2 U7220 ( .A(n4887), .B(n4875), .C(n4809), .Z(n4810) );
  HS65_LH_AOI21X2 U7221 ( .A(n5229), .B(n5658), .C(n4547), .Z(n4567) );
  HS65_LH_NAND2X4 U7222 ( .A(n3634), .B(n5194), .Z(n3636) );
  HS65_LH_IVX9 U7226 ( .A(n5630), .Z(n4419) );
  HS65_LH_NAND3X3 U7227 ( .A(n5563), .B(n5574), .C(n5562), .Z(n5577) );
  HS65_LH_AOI21X2 U7228 ( .A(n5575), .B(n5574), .C(n5573), .Z(n5576) );
  HS65_LH_OAI21X3 U7229 ( .A(n4134), .B(n4795), .C(n4163), .Z(n4381) );
  HS65_LH_AOI21X2 U7230 ( .A(n5304), .B(n5303), .C(n5302), .Z(n5486) );
  HS65_LH_IVX9 U7231 ( .A(n4955), .Z(n4164) );
  HS65_LH_AOI21X2 U7232 ( .A(n4625), .B(n4632), .C(n4627), .Z(n4159) );
  HS65_LH_AOI21X2 U7234 ( .A(n4508), .B(n4943), .C(n4261), .Z(n4260) );
  HS65_LL_OR2X4 U7235 ( .A(n3485), .B(n3484), .Z(n2924) );
  HS65_LL_NAND2AX4 U7236 ( .A(n3246), .B(n3362), .Z(n3894) );
  HS65_LH_IVX4 U7237 ( .A(n4558), .Z(n4157) );
  HS65_LL_OAI12X2 U7238 ( .A(n5046), .B(n5045), .C(n5044), .Z(n5074) );
  HS65_LL_NOR2AX3 U7239 ( .A(n3453), .B(n3452), .Z(n3454) );
  HS65_LH_OAI21X3 U7240 ( .A(n4808), .B(n5656), .C(n4807), .Z(n4809) );
  HS65_LH_AOI21X2 U7241 ( .A(n3704), .B(n5630), .C(n3703), .Z(n3705) );
  HS65_LH_NOR2X5 U7242 ( .A(n4307), .B(n4330), .Z(n4309) );
  HS65_LL_NAND2X2 U7246 ( .A(n4996), .B(n5015), .Z(n5018) );
  HS65_LH_CNIVX3 U7247 ( .A(n3804), .Z(n3685) );
  HS65_LH_AOI21X2 U7248 ( .A(n4424), .B(n5607), .C(n4375), .Z(n4376) );
  HS65_LL_OAI112X1 U7249 ( .A(n5554), .B(n5553), .C(n5552), .D(n5551), .Z(
        n5555) );
  HS65_LH_AOI21X2 U7250 ( .A(n5618), .B(n4892), .C(n4891), .Z(n4893) );
  HS65_LH_AOI21X2 U7251 ( .A(n4943), .B(n4528), .C(n4527), .Z(n4529) );
  HS65_LH_CNIVX3 U7252 ( .A(n5366), .Z(n5291) );
  HS65_LL_NOR2X2 U7253 ( .A(n5646), .B(n5172), .Z(n4434) );
  HS65_LL_AOI21X2 U7254 ( .A(n9352), .B(n5567), .C(n5649), .Z(n3774) );
  HS65_LH_AOI21X2 U7256 ( .A(n9349), .B(n5654), .C(n5649), .Z(n5651) );
  HS65_LH_IVX7 U7257 ( .A(n4872), .Z(n4119) );
  HS65_LH_AND2X4 U7258 ( .A(n3893), .B(n3892), .Z(n2907) );
  HS65_LL_NOR2AX3 U7259 ( .A(n3652), .B(n3651), .Z(n4025) );
  HS65_LH_OAI21X3 U7260 ( .A(n5176), .B(n4800), .C(n4799), .Z(n4815) );
  HS65_LH_AOI21X2 U7261 ( .A(n3921), .B(n3920), .C(n5241), .Z(n3925) );
  HS65_LL_NOR2AX3 U7262 ( .A(n3912), .B(n3911), .Z(n3913) );
  HS65_LH_CNIVX3 U7263 ( .A(n5464), .Z(n5330) );
  HS65_LL_OAI12X2 U7264 ( .A(n5441), .B(n5440), .C(n5439), .Z(n5459) );
  HS65_LH_CNIVX3 U7265 ( .A(n4886), .Z(n4070) );
  HS65_LH_AOI21X2 U7266 ( .A(n5608), .B(n5607), .C(n5606), .Z(n5609) );
  HS65_LL_OAI12X2 U7267 ( .A(n5499), .B(n5346), .C(n5286), .Z(n5575) );
  HS65_LH_AOI21X2 U7268 ( .A(n5234), .B(n3662), .C(n3661), .Z(n3678) );
  HS65_LH_NAND2AX7 U7269 ( .A(n3766), .B(n3765), .Z(n4515) );
  HS65_LH_OAI12X3 U7270 ( .A(n4915), .B(n3891), .C(n3893), .Z(n3367) );
  HS65_LLS_XOR2X3 U7271 ( .A(n9202), .B(n7800), .Z(
        \u_DataPath/u_execute/link_value_i [31]) );
  HS65_LL_NAND3X3 U7272 ( .A(n3821), .B(n3781), .C(n3780), .Z(n5644) );
  HS65_LH_AND2X4 U7273 ( .A(n5435), .B(n5628), .Z(n2917) );
  HS65_LH_NAND2X7 U7274 ( .A(n3499), .B(n5608), .Z(n3501) );
  HS65_LL_OAI12X3 U7276 ( .A(n4257), .B(n4256), .C(n3426), .Z(n4262) );
  HS65_LH_OAI12X3 U7277 ( .A(n4630), .B(n4629), .C(n4628), .Z(n4631) );
  HS65_LH_NAND3X5 U7278 ( .A(n3833), .B(n3832), .C(n3831), .Z(n5142) );
  HS65_LL_NAND2AX4 U7279 ( .A(n3528), .B(n3527), .Z(n4393) );
  HS65_LH_CNIVX3 U7280 ( .A(n4748), .Z(n3919) );
  HS65_LH_NAND2AX4 U7281 ( .A(n3981), .B(n5615), .Z(n3792) );
  HS65_LHS_XOR2X6 U7282 ( .A(n5742), .B(n5854), .Z(\u_DataPath/toPC2_i [30])
         );
  HS65_LL_NOR2AX3 U7283 ( .A(n3197), .B(n4244), .Z(n3374) );
  HS65_LL_NAND2X4 U7284 ( .A(n4724), .B(n5423), .Z(n5346) );
  HS65_LL_AOI22X1 U7286 ( .A(n8868), .B(n9180), .C(n9368), .D(n8869), .Z(n8395) );
  HS65_LL_OAI12X3 U7287 ( .A(n5193), .B(n3572), .C(n3574), .Z(n3750) );
  HS65_LH_AOI31X2 U7288 ( .A(n2854), .B(n5567), .C(n5566), .D(n5565), .Z(n5578) );
  HS65_LL_NAND3X2 U7289 ( .A(n4061), .B(n3664), .C(n3663), .Z(n5228) );
  HS65_LH_OAI12X3 U7290 ( .A(n4038), .B(n4034), .C(n4036), .Z(n3476) );
  HS65_LH_AOI21X2 U7292 ( .A(n4587), .B(n2858), .C(n3957), .Z(n3958) );
  HS65_LH_AOI21X2 U7293 ( .A(n4975), .B(n4974), .C(n5499), .Z(n4996) );
  HS65_LH_NOR2AX3 U7294 ( .A(n3231), .B(n4902), .Z(n4014) );
  HS65_LL_NAND2AX4 U7295 ( .A(n3361), .B(n4904), .Z(n4016) );
  HS65_LL_NOR2X3 U7297 ( .A(\sub_x_53/A[25] ), .B(n5425), .Z(n3572) );
  HS65_LH_AOI21X2 U7298 ( .A(n3426), .B(n4066), .C(n3969), .Z(n4894) );
  HS65_LH_NAND2X4 U7299 ( .A(n3700), .B(n3699), .Z(n3708) );
  HS65_LH_NAND2X4 U7300 ( .A(n4641), .B(n4142), .Z(n4146) );
  HS65_LL_AOI22X1 U7301 ( .A(\sub_x_53/A[25] ), .B(n4551), .C(n2845), .D(
        \lte_x_59/B[24] ), .Z(n3602) );
  HS65_LL_AOI22X1 U7302 ( .A(n8868), .B(n9266), .C(n9365), .D(n8870), .Z(n8445) );
  HS65_LH_NAND2X4 U7303 ( .A(n7631), .B(n5124), .Z(n5157) );
  HS65_LL_NOR2X2 U7304 ( .A(n3731), .B(n5603), .Z(n3499) );
  HS65_LH_AOI21X2 U7305 ( .A(n9352), .B(n4674), .C(n4067), .Z(n4069) );
  HS65_LH_NAND2AX4 U7307 ( .A(n4643), .B(n3330), .Z(n3351) );
  HS65_LL_OAI12X3 U7309 ( .A(n4882), .B(n4876), .C(n4878), .Z(n4040) );
  HS65_LH_AO22X9 U7310 ( .A(n8905), .B(n9188), .C(n9133), .D(n8998), .Z(
        \u_DataPath/jump_address_i [28]) );
  HS65_LL_AOI12X2 U7311 ( .A(n4824), .B(n5126), .C(n4596), .Z(n3487) );
  HS65_LH_NAND2X4 U7312 ( .A(n5258), .B(n5261), .Z(n4253) );
  HS65_LH_AOI31X2 U7313 ( .A(\sub_x_53/A[25] ), .B(n5345), .C(n5344), .D(n5343), .Z(n5349) );
  HS65_LH_AND2X4 U7315 ( .A(n4036), .B(n4035), .Z(n4045) );
  HS65_LH_AOI31X2 U7316 ( .A(\lte_x_59/B[7] ), .B(n5313), .C(n5312), .D(n5311), 
        .Z(n5314) );
  HS65_LH_OAI21X2 U7317 ( .A(n5435), .B(n3698), .C(n5509), .Z(n5436) );
  HS65_LHS_XNOR2X6 U7318 ( .A(n5861), .B(n5860), .Z(\u_DataPath/toPC2_i [29])
         );
  HS65_LL_NOR2X2 U7319 ( .A(n4968), .B(n5361), .Z(n5009) );
  HS65_LH_AOI21X2 U7320 ( .A(n4551), .B(\lte_x_59/B[15] ), .C(n3907), .Z(n3912) );
  HS65_LH_OAI21X3 U7321 ( .A(n5318), .B(n5037), .C(n5317), .Z(n5554) );
  HS65_LHS_XNOR2X6 U7323 ( .A(n6056), .B(n6055), .Z(
        \u_DataPath/u_execute/resAdd1_i [30]) );
  HS65_LH_OAI21X2 U7324 ( .A(n5065), .B(n5064), .C(n5063), .Z(n5066) );
  HS65_LH_AOI21X2 U7325 ( .A(n4551), .B(\sub_x_53/A[25] ), .C(n3549), .Z(n3585) );
  HS65_LH_OAI22X3 U7326 ( .A(n7306), .B(n8337), .C(n7915), .D(n8336), .Z(
        \u_DataPath/data_read_ex_1_i [9]) );
  HS65_LH_OAI22X3 U7327 ( .A(n7306), .B(n8330), .C(n7915), .D(n8329), .Z(
        \u_DataPath/data_read_ex_1_i [25]) );
  HS65_LH_OAI22X3 U7328 ( .A(n7306), .B(n8444), .C(n7914), .D(n8173), .Z(
        \u_DataPath/data_read_ex_1_i [2]) );
  HS65_LH_AND2X4 U7329 ( .A(\lte_x_59/B[9] ), .B(n2864), .Z(n4153) );
  HS65_LH_AO22X9 U7330 ( .A(n9255), .B(n9188), .C(n9133), .D(n9013), .Z(
        \u_DataPath/jump_address_i [9]) );
  HS65_LH_AO222X4 U7331 ( .A(\u_DataPath/pc_4_i [31]), .B(n7896), .C(n7887), 
        .D(n9165), .E(n7893), .F(n9403), .Z(n8641) );
  HS65_LH_OAI22X3 U7334 ( .A(n4981), .B(n5129), .C(n2854), .D(n3756), .Z(n3782) );
  HS65_LL_OAI12X3 U7335 ( .A(n4418), .B(n4407), .C(n5434), .Z(n5629) );
  HS65_LH_OR2X4 U7336 ( .A(\sub_x_53/A[0] ), .B(n5136), .Z(n5125) );
  HS65_LH_NAND3X2 U7337 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5531), .C(n5506), 
        .Z(n5080) );
  HS65_LH_NOR2X5 U7338 ( .A(n2858), .B(n5398), .Z(n5399) );
  HS65_LL_NOR2X2 U7339 ( .A(n5430), .B(n4244), .Z(n5432) );
  HS65_LL_NOR2X3 U7340 ( .A(n5419), .B(n4407), .Z(n5632) );
  HS65_LL_OR2X4 U7341 ( .A(n5021), .B(n5022), .Z(n2892) );
  HS65_LH_NOR2AX3 U7343 ( .A(n4682), .B(n3360), .Z(n4905) );
  HS65_LL_NOR2X3 U7344 ( .A(n2843), .B(n4683), .Z(n5300) );
  HS65_LH_NOR2X5 U7345 ( .A(n4676), .B(n5061), .Z(n5083) );
  HS65_LH_NAND2X5 U7346 ( .A(n5031), .B(n5030), .Z(n5544) );
  HS65_LH_NOR2X3 U7347 ( .A(n5320), .B(n5321), .Z(n5037) );
  HS65_LH_NOR2X5 U7348 ( .A(n4811), .B(n4805), .Z(n5548) );
  HS65_LH_NOR2X5 U7349 ( .A(n5031), .B(n5030), .Z(n5095) );
  HS65_LH_NAND2X5 U7350 ( .A(n3101), .B(n4997), .Z(n5289) );
  HS65_LH_NOR2X5 U7351 ( .A(n4711), .B(n4976), .Z(n5347) );
  HS65_LL_NOR2X2 U7352 ( .A(n4701), .B(n5418), .Z(n5363) );
  HS65_LH_NOR2AX3 U7353 ( .A(n5004), .B(n3372), .Z(n5269) );
  HS65_LH_OAI12X3 U7354 ( .A(n4628), .B(n4622), .C(n4624), .Z(n3485) );
  HS65_LL_NAND2X4 U7355 ( .A(\sub_x_53/A[0] ), .B(n5136), .Z(n5126) );
  HS65_LH_NOR4ABX2 U7357 ( .A(n7406), .B(n7405), .C(n7404), .D(n7403), .Z(
        n8433) );
  HS65_LH_NOR4ABX2 U7358 ( .A(n7471), .B(n7470), .C(n7469), .D(n7468), .Z(
        n8373) );
  HS65_LH_NOR4ABX2 U7359 ( .A(n7386), .B(n7385), .C(n7384), .D(n7383), .Z(
        n8388) );
  HS65_LH_NOR4ABX2 U7360 ( .A(n7451), .B(n7450), .C(n7449), .D(n7448), .Z(
        n8155) );
  HS65_LH_NOR4ABX2 U7361 ( .A(n7557), .B(n7556), .C(n7555), .D(n7554), .Z(
        n8354) );
  HS65_LH_NOR4ABX2 U7362 ( .A(n7612), .B(n7611), .C(n7610), .D(n7609), .Z(
        n8363) );
  HS65_LH_NOR4ABX2 U7363 ( .A(n6204), .B(n6203), .C(n6202), .D(n6201), .Z(
        n8366) );
  HS65_LH_NOR4ABX2 U7364 ( .A(n6494), .B(n6493), .C(n6492), .D(n6491), .Z(
        n8313) );
  HS65_LH_NOR4ABX2 U7365 ( .A(n6325), .B(n6324), .C(n6323), .D(n6322), .Z(
        n8403) );
  HS65_LH_NOR4ABX2 U7366 ( .A(n7366), .B(n7365), .C(n7364), .D(n7363), .Z(
        n8392) );
  HS65_LH_NOR4ABX2 U7367 ( .A(n7537), .B(n7536), .C(n7535), .D(n7534), .Z(
        n8381) );
  HS65_LH_NOR4ABX2 U7368 ( .A(n7577), .B(n7576), .C(n7575), .D(n7574), .Z(
        n8368) );
  HS65_LH_NOR4ABX2 U7369 ( .A(n6975), .B(n6974), .C(n6973), .D(n6972), .Z(
        n8442) );
  HS65_LH_NOR4ABX2 U7370 ( .A(n6304), .B(n6303), .C(n6302), .D(n6301), .Z(
        n8371) );
  HS65_LH_NOR4ABX2 U7371 ( .A(n7491), .B(n7490), .C(n7489), .D(n7488), .Z(
        n8384) );
  HS65_LH_NOR4ABX2 U7372 ( .A(n6161), .B(n6160), .C(n6159), .D(n6158), .Z(
        n8396) );
  HS65_LH_NOR4ABX2 U7373 ( .A(n6284), .B(n6283), .C(n6282), .D(n6281), .Z(
        n8352) );
  HS65_LH_NOR4ABX2 U7374 ( .A(n7427), .B(n7426), .C(n7425), .D(n7424), .Z(
        n8379) );
  HS65_LH_NOR4ABX2 U7375 ( .A(n7511), .B(n7510), .C(n7509), .D(n7508), .Z(
        n8382) );
  HS65_LH_AO22X9 U7377 ( .A(n8997), .B(n9188), .C(n9133), .D(n9011), .Z(
        \u_DataPath/jump_address_i [7]) );
  HS65_LH_OR2X4 U7380 ( .A(n2851), .B(n7623), .Z(n4205) );
  HS65_LH_AO22X9 U7382 ( .A(n9022), .B(n9188), .C(n9133), .D(n8948), .Z(
        \u_DataPath/jump_address_i [14]) );
  HS65_LH_NOR2X5 U7383 ( .A(\sub_x_53/A[2] ), .B(n5088), .Z(n4596) );
  HS65_LH_AO22X9 U7384 ( .A(n9055), .B(n9188), .C(n9133), .D(n8934), .Z(
        \u_DataPath/jump_address_i [24]) );
  HS65_LH_AO22X9 U7388 ( .A(n9260), .B(n9188), .C(n9133), .D(n9054), .Z(
        \u_DataPath/jump_address_i [26]) );
  HS65_LH_AO222X4 U7389 ( .A(n7896), .B(\u_DataPath/pc_4_i [30]), .C(n7893), 
        .D(\u_DataPath/jump_address_i [30]), .E(n9025), .F(n7887), .Z(n8642)
         );
  HS65_LH_IVX9 U7390 ( .A(n4550), .Z(n4863) );
  HS65_LL_NOR2X3 U7391 ( .A(n4726), .B(n4966), .Z(n5503) );
  HS65_LH_IVX9 U7392 ( .A(\lte_x_59/B[4] ), .Z(n4796) );
  HS65_LH_AOI21X2 U7400 ( .A(n5648), .B(n4147), .C(n5647), .Z(n4165) );
  HS65_LH_IVX9 U7402 ( .A(n4458), .Z(n4949) );
  HS65_LL_NOR2AX6 U7403 ( .A(n5088), .B(n3425), .Z(n3426) );
  HS65_LH_NOR2X6 U7406 ( .A(n7785), .B(n7784), .Z(n7786) );
  HS65_LL_OAI12X3 U7407 ( .A(n5952), .B(n5955), .C(n5954), .Z(n6119) );
  HS65_LH_OAI21X3 U7410 ( .A(n9246), .B(n8453), .C(n9086), .Z(
        \u_DataPath/from_mem_data_out_i [28]) );
  HS65_LL_NOR2X6 U7416 ( .A(n3106), .B(n3105), .Z(\lte_x_59/B[7] ) );
  HS65_LH_IVX9 U7417 ( .A(n4699), .Z(n3376) );
  HS65_LL_AO12X4 U7418 ( .A(n3274), .B(n3270), .C(n3269), .Z(n2925) );
  HS65_LH_IVX9 U7419 ( .A(n4967), .Z(n5417) );
  HS65_LH_AO222X4 U7420 ( .A(n7896), .B(\u_DataPath/pc_4_i [24]), .C(n7893), 
        .D(\u_DataPath/jump_address_i [24]), .E(n8931), .F(n7887), .Z(n8648)
         );
  HS65_LHS_XOR2X3 U7421 ( .A(n7795), .B(n7794), .Z(
        \u_DataPath/u_execute/link_value_i [27]) );
  HS65_LH_AO222X4 U7422 ( .A(n7896), .B(\u_DataPath/pc_4_i [29]), .C(n7893), 
        .D(n9417), .E(n9164), .F(n7887), .Z(n8643) );
  HS65_LH_AO222X4 U7423 ( .A(n7895), .B(\u_DataPath/pc_4_i [17]), .C(n7892), 
        .D(n9406), .E(n8928), .F(n7888), .Z(n8655) );
  HS65_LH_IVX9 U7424 ( .A(n5021), .Z(n4985) );
  HS65_LH_AO22X9 U7425 ( .A(n9254), .B(n8797), .C(n9240), .D(n8992), .Z(
        \u_DataPath/pc4_to_idexreg_i [24]) );
  HS65_LH_AO22X9 U7426 ( .A(n9254), .B(n8796), .C(n9132), .D(n8993), .Z(
        \u_DataPath/pc4_to_idexreg_i [29]) );
  HS65_LH_AO22X9 U7427 ( .A(n9254), .B(n8795), .C(n9240), .D(n8994), .Z(
        \u_DataPath/pc4_to_idexreg_i [17]) );
  HS65_LL_NAND2AX7 U7428 ( .A(n2922), .B(n3277), .Z(n5062) );
  HS65_LH_AOI22X3 U7430 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][18] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][18] ), .Z(n6344)
         );
  HS65_LH_OAI22X6 U7431 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [21]), .C(
        n8364), .D(n3409), .Z(n3060) );
  HS65_LL_NAND2X5 U7432 ( .A(n3164), .B(n3163), .Z(n4967) );
  HS65_LH_IVX9 U7433 ( .A(n5654), .Z(n2869) );
  HS65_LH_NOR2X5 U7434 ( .A(n9399), .B(n3341), .Z(n3066) );
  HS65_LH_AO22X9 U7435 ( .A(n8793), .B(n9138), .C(n9331), .D(n9153), .Z(
        opcode_i[3]) );
  HS65_LH_AO22X9 U7436 ( .A(n8792), .B(n9138), .C(n9329), .D(n9153), .Z(
        opcode_i[1]) );
  HS65_LH_NAND2X4 U7437 ( .A(n9281), .B(n8399), .Z(n8273) );
  HS65_LH_NAND2X4 U7438 ( .A(n9282), .B(n8399), .Z(n8334) );
  HS65_LH_AO22X9 U7439 ( .A(n8791), .B(n9252), .C(n9317), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [14]) );
  HS65_LH_NAND2X4 U7440 ( .A(n9283), .B(n8399), .Z(n8295) );
  HS65_LH_AO22X9 U7441 ( .A(n8790), .B(n9252), .C(n9316), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [13]) );
  HS65_LH_NAND2X4 U7442 ( .A(n9284), .B(n8399), .Z(n8346) );
  HS65_LH_AO22X9 U7443 ( .A(n8789), .B(n9252), .C(n9315), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [12]) );
  HS65_LH_AO22X9 U7444 ( .A(n8788), .B(n9252), .C(n9314), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [11]) );
  HS65_LH_NAND2X4 U7446 ( .A(n9286), .B(n8399), .Z(n8341) );
  HS65_LH_NAND2X4 U7447 ( .A(n9287), .B(n8399), .Z(n8400) );
  HS65_LH_NAND2X4 U7448 ( .A(n9288), .B(n8399), .Z(n8308) );
  HS65_LH_AO22X9 U7449 ( .A(n8787), .B(n9252), .C(n9321), .D(n9141), .Z(
        \u_DataPath/jaddr_i [18]) );
  HS65_LH_BFX9 U7451 ( .A(n8443), .Z(n7901) );
  HS65_LHS_XNOR2X6 U7452 ( .A(n7705), .B(n7780), .Z(\u_DataPath/pc_4_i [29])
         );
  HS65_LH_AO222X4 U7453 ( .A(n7895), .B(\u_DataPath/pc_4_i [22]), .C(n7892), 
        .D(\u_DataPath/jump_address_i [22]), .E(n8929), .F(n7887), .Z(n8650)
         );
  HS65_LL_OR2X4 U7455 ( .A(n8800), .B(n3341), .Z(n2903) );
  HS65_LH_AO222X4 U7457 ( .A(n7896), .B(\u_DataPath/pc_4_i [28]), .C(n7893), 
        .D(\u_DataPath/jump_address_i [28]), .E(n8941), .F(n7887), .Z(n8644)
         );
  HS65_LH_OAI22X6 U7458 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [12]), .C(
        n8255), .D(n3409), .Z(n3265) );
  HS65_LL_NAND2X5 U7459 ( .A(n3263), .B(n3262), .Z(n5048) );
  HS65_LH_AO22X9 U7460 ( .A(n8785), .B(n9138), .C(n9322), .D(n9153), .Z(
        \u_DataPath/jaddr_i [19]) );
  HS65_LH_AO22X9 U7462 ( .A(n8784), .B(n9253), .C(n9310), .D(n9142), .Z(
        \u_DataPath/immediate_ext_dec_i [7]) );
  HS65_LH_AO22X9 U7463 ( .A(n8783), .B(n9253), .C(n9311), .D(n9142), .Z(
        \u_DataPath/immediate_ext_dec_i [8]) );
  HS65_LH_AO22X9 U7465 ( .A(n8781), .B(n9253), .C(n9313), .D(n9142), .Z(
        \u_DataPath/immediate_ext_dec_i [10]) );
  HS65_LH_AO22X9 U7467 ( .A(n8779), .B(n9252), .C(n9308), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [5]) );
  HS65_LH_AO22X9 U7468 ( .A(n8778), .B(n9252), .C(n9309), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [6]) );
  HS65_LH_AO222X4 U7469 ( .A(n7895), .B(\u_DataPath/pc_4_i [23]), .C(n7892), 
        .D(n9414), .E(n9197), .F(n7887), .Z(n8649) );
  HS65_LH_NAND2X7 U7470 ( .A(n9207), .B(n7122), .Z(n7794) );
  HS65_LH_AO222X4 U7471 ( .A(n7895), .B(\u_DataPath/pc_4_i [21]), .C(n7892), 
        .D(n9405), .E(n9193), .F(n7887), .Z(n8651) );
  HS65_LH_AO222X4 U7472 ( .A(n7895), .B(\u_DataPath/pc_4_i [16]), .C(n7892), 
        .D(\u_DataPath/jump_address_i [16]), .E(n9194), .F(n7888), .Z(n8656)
         );
  HS65_LHS_XNOR2X6 U7474 ( .A(n3121), .B(n7687), .Z(\u_DataPath/pc_4_i [24])
         );
  HS65_LH_AO22X9 U7475 ( .A(n8776), .B(n9252), .C(n9303), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [0]) );
  HS65_LH_AO22X9 U7477 ( .A(n8772), .B(n9252), .C(n9306), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [3]) );
  HS65_LHS_XOR2X6 U7479 ( .A(n7769), .B(n7768), .Z(\u_DataPath/pc_4_i [21]) );
  HS65_LHS_XOR2X3 U7481 ( .A(n5975), .B(n5974), .Z(
        \u_DataPath/u_execute/resAdd1_i [25]) );
  HS65_LH_OAI21X3 U7482 ( .A(n8494), .B(n8390), .C(n8493), .Z(
        \u_DataPath/mem_writedata_out_i [4]) );
  HS65_LHS_XOR2X6 U7483 ( .A(n7766), .B(n7765), .Z(\u_DataPath/pc_4_i [23]) );
  HS65_LL_AO12X4 U7484 ( .A(n3414), .B(n8491), .C(n3413), .Z(n3425) );
  HS65_LL_NAND3AX3 U7485 ( .A(n3162), .B(n3161), .C(n8548), .Z(n3163) );
  HS65_LHS_XOR2X6 U7486 ( .A(n7756), .B(n7755), .Z(\u_DataPath/pc_4_i [22]) );
  HS65_LHS_XOR2X3 U7487 ( .A(n7799), .B(n7798), .Z(
        \u_DataPath/u_execute/link_value_i [25]) );
  HS65_LL_OR2X4 U7488 ( .A(n3171), .B(n8544), .Z(n2905) );
  HS65_LH_AO222X4 U7489 ( .A(n7896), .B(\u_DataPath/pc_4_i [27]), .C(n7893), 
        .D(n9416), .E(n9264), .F(n7887), .Z(n8645) );
  HS65_LH_BFX9 U7490 ( .A(n8482), .Z(n7920) );
  HS65_LH_NOR3X2 U7491 ( .A(n8773), .B(n9099), .C(n8114), .Z(n8129) );
  HS65_LH_NOR2X3 U7492 ( .A(n9083), .B(n8916), .Z(\u_DataPath/cw_exmem_i [6])
         );
  HS65_LHS_XOR2X6 U7493 ( .A(n3122), .B(n7754), .Z(\u_DataPath/pc_4_i [16]) );
  HS65_LL_NOR3X1 U7495 ( .A(n8775), .B(n9169), .C(n8114), .Z(n8082) );
  HS65_LL_NOR3X1 U7496 ( .A(n8771), .B(n9003), .C(n8114), .Z(n8106) );
  HS65_LL_NAND3X3 U7497 ( .A(n4714), .B(n8562), .C(n8561), .Z(n4974) );
  HS65_LL_OA31X4 U7498 ( .A(n9401), .B(n3288), .C(n4713), .D(n3287), .Z(n2910)
         );
  HS65_LL_NAND2AX4 U7499 ( .A(n3194), .B(n8532), .Z(n3196) );
  HS65_LL_NAND3AX3 U7501 ( .A(n3228), .B(n3227), .C(n6124), .Z(n3229) );
  HS65_LL_OAI22X3 U7502 ( .A(n3333), .B(\u_DataPath/dataOut_exe_i [6]), .C(
        n8311), .D(n3340), .Z(n3319) );
  HS65_LHS_XNOR2X6 U7503 ( .A(n2831), .B(n7767), .Z(\u_DataPath/pc_4_i [20])
         );
  HS65_LHS_XNOR2X6 U7504 ( .A(n3123), .B(n7677), .Z(\u_DataPath/pc_4_i [14])
         );
  HS65_LHS_XNOR2X3 U7505 ( .A(n7121), .B(n7120), .Z(
        \u_DataPath/u_execute/link_value_i [24]) );
  HS65_LH_NAND2X7 U7506 ( .A(n3292), .B(n3291), .Z(n3397) );
  HS65_LHS_XNOR2X6 U7507 ( .A(n6068), .B(n6067), .Z(
        \u_DataPath/u_execute/resAdd1_i [19]) );
  HS65_LL_OAI22X3 U7508 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [8]), .C(
        n8265), .D(n3340), .Z(n3213) );
  HS65_LL_OAI12X12 U7509 ( .A(n8141), .B(n8147), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N151 ) );
  HS65_LH_NAND2X5 U7510 ( .A(n2896), .B(n3189), .Z(n8534) );
  HS65_LHS_XNOR2X6 U7511 ( .A(n9357), .B(n7655), .Z(\u_DataPath/pc_4_i [13])
         );
  HS65_LL_OAI13X5 U7512 ( .A(n3329), .B(n8501), .C(n8500), .D(n3328), .Z(n5030) );
  HS65_LH_AND2X4 U7513 ( .A(n4714), .B(n8521), .Z(n3279) );
  HS65_LL_OAI12X18 U7514 ( .A(n8147), .B(n8150), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N135 ) );
  HS65_LH_NAND2X4 U7515 ( .A(n8566), .B(n8484), .Z(n7870) );
  HS65_LL_OAI12X12 U7516 ( .A(n8145), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N125 ) );
  HS65_LL_OAI12X18 U7517 ( .A(n3009), .B(n8150), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N132 ) );
  HS65_LH_BFX9 U7518 ( .A(n8456), .Z(n7914) );
  HS65_LL_OAI12X18 U7519 ( .A(n3010), .B(n8150), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N137 ) );
  HS65_LH_NAND3X3 U7520 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .B(n8120), 
        .C(n8635), .Z(n8077) );
  HS65_LH_AOI12X2 U7521 ( .A(n6057), .B(n6059), .C(n5764), .Z(n5969) );
  HS65_LHS_XNOR2X6 U7522 ( .A(n3120), .B(n7674), .Z(\u_DataPath/pc_4_i [25])
         );
  HS65_LL_NAND2AX4 U7523 ( .A(n7878), .B(n4212), .Z(n4216) );
  HS65_LL_NOR3X1 U7525 ( .A(n8542), .B(n4713), .C(n8541), .Z(n3181) );
  HS65_LH_BFX9 U7526 ( .A(n8456), .Z(n7916) );
  HS65_LH_BFX9 U7527 ( .A(n8456), .Z(n7915) );
  HS65_LL_OAI12X12 U7528 ( .A(n3012), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N126 ) );
  HS65_LL_NOR4ABX2 U7529 ( .A(n8269), .B(n8318), .C(n9235), .D(n8268), .Z(
        n8272) );
  HS65_LH_OAI21X3 U7530 ( .A(n8098), .B(n8097), .C(n8635), .Z(n8094) );
  HS65_LL_NOR2AX3 U7532 ( .A(n3219), .B(n3218), .Z(n5693) );
  HS65_LH_BFX9 U7533 ( .A(n8287), .Z(n7896) );
  HS65_LH_BFX9 U7535 ( .A(n8287), .Z(n7894) );
  HS65_LL_OAI21X2 U7536 ( .A(n3284), .B(n4714), .C(n3283), .Z(n3289) );
  HS65_LH_OAI12X3 U7537 ( .A(n5763), .B(n5773), .C(n5762), .Z(n5864) );
  HS65_LL_NAND2X7 U7538 ( .A(n7306), .B(n7095), .Z(n7096) );
  HS65_LH_OAI12X3 U7539 ( .A(n6066), .B(n6065), .C(n6064), .Z(n6067) );
  HS65_LHS_XOR2X3 U7540 ( .A(n6030), .B(n6029), .Z(
        \u_DataPath/u_execute/resAdd1_i [23]) );
  HS65_LH_BFX9 U7541 ( .A(n8287), .Z(n7895) );
  HS65_LH_AND2X4 U7542 ( .A(n8537), .B(n2866), .Z(n2894) );
  HS65_LL_OAI12X3 U7543 ( .A(n6026), .B(n6029), .C(n6028), .Z(n6107) );
  HS65_LL_NAND2AX4 U7544 ( .A(n8332), .B(n2866), .Z(n8505) );
  HS65_LL_OA12X4 U7545 ( .A(n4713), .B(n3347), .C(n3346), .Z(n3348) );
  HS65_LHS_XOR2X3 U7546 ( .A(n3119), .B(n7759), .Z(\u_DataPath/pc_4_i [26]) );
  HS65_LH_BFX9 U7547 ( .A(n8483), .Z(n7924) );
  HS65_LHS_XOR2X3 U7548 ( .A(n7797), .B(n7796), .Z(
        \u_DataPath/u_execute/link_value_i [23]) );
  HS65_LH_NOR2X3 U7549 ( .A(n8719), .B(n4712), .Z(n7878) );
  HS65_LL_NAND3X3 U7550 ( .A(n8143), .B(n7619), .C(n7618), .Z(n8148) );
  HS65_LH_NOR2X5 U7552 ( .A(n8716), .B(n7802), .Z(n3299) );
  HS65_LH_IVX9 U7553 ( .A(n7661), .Z(n7757) );
  HS65_LL_AOI12X6 U7554 ( .A(n8161), .B(n8160), .C(n8159), .Z(
        \u_DataPath/u_idexreg/N184 ) );
  HS65_LH_NAND2X4 U7556 ( .A(n8297), .B(n7802), .Z(n8502) );
  HS65_LH_NAND2X7 U7557 ( .A(n3110), .B(n8132), .Z(n8573) );
  HS65_LH_NAND2X4 U7559 ( .A(n4187), .B(n7802), .Z(n8572) );
  HS65_LH_NOR2X5 U7560 ( .A(n8176), .B(n9401), .Z(n8570) );
  HS65_LH_AOI12X2 U7561 ( .A(n5814), .B(n5868), .C(n5813), .Z(n5815) );
  HS65_LH_NAND2X4 U7562 ( .A(n8681), .B(n7749), .Z(n7750) );
  HS65_LH_NOR2X3 U7563 ( .A(n8364), .B(n9401), .Z(n8542) );
  HS65_LH_NOR2X3 U7564 ( .A(n8350), .B(n9401), .Z(n8544) );
  HS65_LH_AOI12X2 U7565 ( .A(n6005), .B(n5791), .C(n5790), .Z(n5793) );
  HS65_LH_NAND2X5 U7566 ( .A(n3225), .B(n7802), .Z(n8506) );
  HS65_LH_OR2X4 U7567 ( .A(n8426), .B(n9401), .Z(n4212) );
  HS65_LH_AOI12X2 U7569 ( .A(n6069), .B(n5872), .C(n5984), .Z(n5784) );
  HS65_LHS_XNOR2X6 U7570 ( .A(n5889), .B(n5888), .Z(\u_DataPath/toPC2_i [7])
         );
  HS65_LH_NOR2X3 U7571 ( .A(n8374), .B(n9401), .Z(n8559) );
  HS65_LH_AOI12X2 U7572 ( .A(n6005), .B(n5992), .C(n5790), .Z(n5993) );
  HS65_LH_AOI31X3 U7573 ( .A(n9117), .B(n9334), .C(n8714), .D(n8424), .Z(n7847) );
  HS65_LH_OAI12X3 U7574 ( .A(n5887), .B(n5886), .C(n5885), .Z(n5888) );
  HS65_LH_IVX9 U7576 ( .A(n8425), .Z(n8132) );
  HS65_LL_NAND2X2 U7578 ( .A(n3217), .B(n3216), .Z(n3218) );
  HS65_LL_NOR4ABX2 U7579 ( .A(n3053), .B(n3052), .C(n3051), .D(n3034), .Z(
        n3055) );
  HS65_LL_NAND2X7 U7581 ( .A(n8566), .B(n2877), .Z(n8235) );
  HS65_LHS_XOR2X3 U7582 ( .A(n5700), .B(n7710), .Z(n4288) );
  HS65_LH_NAND2X4 U7585 ( .A(n9214), .B(n7729), .Z(n4004) );
  HS65_LH_BFX9 U7586 ( .A(n7886), .Z(n7887) );
  HS65_LH_AOI12X2 U7587 ( .A(n5834), .B(n5892), .C(n5833), .Z(n5886) );
  HS65_LH_BFX9 U7588 ( .A(n7886), .Z(n7888) );
  HS65_LH_AOI31X2 U7589 ( .A(opcode_i[1]), .B(n9084), .C(n7771), .D(n7309), 
        .Z(n8119) );
  HS65_LH_AOI12X2 U7590 ( .A(n6036), .B(n6095), .C(n6035), .Z(n6089) );
  HS65_LH_BFX9 U7592 ( .A(n6683), .Z(n7593) );
  HS65_LH_BFX9 U7593 ( .A(n7886), .Z(n7889) );
  HS65_LH_BFX9 U7594 ( .A(n6746), .Z(n7516) );
  HS65_LH_BFX9 U7595 ( .A(n6172), .Z(n7171) );
  HS65_LH_IVX9 U7596 ( .A(n7861), .Z(n8168) );
  HS65_LH_BFX9 U7597 ( .A(n6754), .Z(n7525) );
  HS65_LH_BFX9 U7600 ( .A(n6635), .Z(n7282) );
  HS65_LH_BFX9 U7602 ( .A(n6680), .Z(n7522) );
  HS65_LH_BFX9 U7603 ( .A(n6171), .Z(n7285) );
  HS65_LH_BFX9 U7607 ( .A(n6739), .Z(n7428) );
  HS65_LH_BFX9 U7608 ( .A(n6634), .Z(n7283) );
  HS65_LH_BFX9 U7609 ( .A(n8285), .Z(n7886) );
  HS65_LL_NOR2X5 U7610 ( .A(n6353), .B(n6333), .Z(n6952) );
  HS65_LL_OAI21X2 U7611 ( .A(n5932), .B(n5963), .C(n5931), .Z(n5933) );
  HS65_LH_BFX9 U7612 ( .A(n7578), .Z(n7429) );
  HS65_LH_BFX9 U7613 ( .A(n6689), .Z(n7603) );
  HS65_LHS_XOR2X6 U7614 ( .A(n7745), .B(n7744), .Z(\u_DataPath/pc_4_i [5]) );
  HS65_LH_BFX9 U7615 ( .A(n6364), .Z(n6927) );
  HS65_LH_OAI211X3 U7617 ( .A(n8089), .B(n7702), .C(n7701), .D(n7700), .Z(
        n8125) );
  HS65_LH_BFX9 U7618 ( .A(n6745), .Z(n7434) );
  HS65_LH_BFX9 U7619 ( .A(n6627), .Z(n7274) );
  HS65_LH_BFX9 U7620 ( .A(n7296), .Z(n6942) );
  HS65_LH_BFX9 U7621 ( .A(n6625), .Z(n7272) );
  HS65_LH_BFX9 U7622 ( .A(n6376), .Z(n7286) );
  HS65_LH_IVX9 U7624 ( .A(n7639), .Z(n7640) );
  HS65_LH_OAI12X3 U7625 ( .A(n5795), .B(n5800), .C(n5797), .Z(n5807) );
  HS65_LL_CB4I1X4 U7626 ( .A(n7834), .B(n5491), .C(n3421), .D(n3422), .Z(n3443) );
  HS65_LHS_XOR2X3 U7627 ( .A(\u_DataPath/jaddr_i [16]), .B(n7089), .Z(n7091)
         );
  HS65_LH_BFX9 U7628 ( .A(n6636), .Z(n7170) );
  HS65_LH_BFX9 U7629 ( .A(n6385), .Z(n7297) );
  HS65_LH_CBI4I1X5 U7630 ( .A(n9084), .B(n7697), .C(n7688), .D(n8084), .Z(
        n7637) );
  HS65_LH_IVX4 U7631 ( .A(n5800), .Z(n5801) );
  HS65_LH_CNIVX3 U7632 ( .A(n7906), .Z(n7849) );
  HS65_LH_BFX9 U7633 ( .A(n6966), .Z(n7333) );
  HS65_LHS_XOR2X6 U7634 ( .A(n8163), .B(n7089), .Z(n7077) );
  HS65_LH_BFX9 U7635 ( .A(n6967), .Z(n7334) );
  HS65_LH_NOR2X2 U7636 ( .A(n9233), .B(n7117), .Z(n7879) );
  HS65_LH_BFX9 U7637 ( .A(n6951), .Z(n7415) );
  HS65_LH_BFX9 U7638 ( .A(n8282), .Z(n7881) );
  HS65_LH_BFX9 U7639 ( .A(n8451), .Z(n7908) );
  HS65_LH_NAND2X4 U7640 ( .A(n5863), .B(n6057), .Z(n5865) );
  HS65_LH_IVX4 U7641 ( .A(n5780), .Z(n5781) );
  HS65_LH_NAND2X4 U7642 ( .A(n6058), .B(n6057), .Z(n6060) );
  HS65_LL_NOR2X5 U7643 ( .A(n6148), .B(n6133), .Z(n6629) );
  HS65_LH_NAND2X4 U7645 ( .A(n6064), .B(n6009), .Z(n6012) );
  HS65_LH_NAND2X4 U7646 ( .A(n6040), .B(n5837), .Z(n6044) );
  HS65_LLS_XNOR2X3 U7647 ( .A(n7618), .B(n3031), .Z(n3054) );
  HS65_LH_NAND2X4 U7648 ( .A(n5876), .B(n5875), .Z(n5881) );
  HS65_LH_NAND2X4 U7649 ( .A(n8685), .B(n7743), .Z(n7744) );
  HS65_LH_BFX9 U7650 ( .A(n7890), .Z(n7891) );
  HS65_LH_BFX9 U7652 ( .A(n7890), .Z(n7893) );
  HS65_LH_NAND2X4 U7653 ( .A(n5896), .B(n6098), .Z(n5901) );
  HS65_LH_NAND2X4 U7654 ( .A(n5848), .B(n6046), .Z(n5849) );
  HS65_LL_NOR2X5 U7655 ( .A(n6153), .B(n6133), .Z(n6370) );
  HS65_LHS_XNOR2X6 U7656 ( .A(n8166), .B(n7618), .Z(n7079) );
  HS65_LH_NAND2X4 U7657 ( .A(n5897), .B(n6050), .Z(n5845) );
  HS65_LH_NAND2X4 U7658 ( .A(n5789), .B(n6005), .Z(n5774) );
  HS65_LL_NOR2X5 U7659 ( .A(n2885), .B(n6133), .Z(n6371) );
  HS65_LH_NAND2X4 U7661 ( .A(n6070), .B(n6069), .Z(n6072) );
  HS65_LL_NOR2X5 U7662 ( .A(n2886), .B(n6132), .Z(n6627) );
  HS65_LH_IVX7 U7664 ( .A(n5121), .Z(n4787) );
  HS65_LH_CNIVX3 U7665 ( .A(n8350), .Z(n3167) );
  HS65_LH_NAND2X4 U7666 ( .A(n5871), .B(n6069), .Z(n5873) );
  HS65_LH_OR2X9 U7667 ( .A(n3345), .B(n4713), .Z(n3349) );
  HS65_LL_NOR2X5 U7668 ( .A(n2885), .B(n6151), .Z(n6364) );
  HS65_LH_AND2X4 U7669 ( .A(n3327), .B(n9183), .Z(n2921) );
  HS65_LL_NAND2AX4 U7670 ( .A(n7619), .B(n2943), .Z(n2945) );
  HS65_LH_CNIVX3 U7671 ( .A(n8550), .Z(n3142) );
  HS65_LH_NAND2X4 U7672 ( .A(n5978), .B(n5977), .Z(n5986) );
  HS65_LH_NAND2X4 U7673 ( .A(n5797), .B(n5796), .Z(n5804) );
  HS65_LH_NAND2X4 U7674 ( .A(n5997), .B(n5996), .Z(n6004) );
  HS65_LH_NAND2X4 U7678 ( .A(n9219), .B(n7789), .Z(n7790) );
  HS65_LH_IVX4 U7679 ( .A(n5981), .Z(n5982) );
  HS65_LH_NAND2X4 U7680 ( .A(n5838), .B(n5837), .Z(n5842) );
  HS65_LH_NAND2X4 U7681 ( .A(n6006), .B(n6005), .Z(n6008) );
  HS65_LH_NAND2X4 U7682 ( .A(n6088), .B(n5831), .Z(n6037) );
  HS65_LL_NOR2X5 U7683 ( .A(n6148), .B(n6147), .Z(n6383) );
  HS65_LH_NAND2X4 U7684 ( .A(n5891), .B(n5890), .Z(n5893) );
  HS65_LH_NAND2X4 U7685 ( .A(n6021), .B(n6020), .Z(n6025) );
  HS65_LLS_XNOR2X3 U7687 ( .A(n9004), .B(n7619), .Z(n3050) );
  HS65_LH_NAND3X3 U7688 ( .A(n8096), .B(n8157), .C(n8076), .Z(n7700) );
  HS65_LL_AND2X4 U7690 ( .A(n2949), .B(n2948), .Z(n2952) );
  HS65_LH_NAND2X4 U7691 ( .A(n6087), .B(n5883), .Z(n6092) );
  HS65_LH_NAND2X4 U7692 ( .A(n5755), .B(n5958), .Z(n5766) );
  HS65_LH_BFX9 U7693 ( .A(n7890), .Z(n7892) );
  HS65_LLS_XNOR2X3 U7694 ( .A(\u_DataPath/jaddr_i [19]), .B(n7619), .Z(n7090)
         );
  HS65_LLS_XNOR2X3 U7695 ( .A(n3029), .B(n7086), .Z(n3048) );
  HS65_LH_NAND2X4 U7696 ( .A(n5745), .B(n5744), .Z(n5747) );
  HS65_LL_NAND2AX7 U7698 ( .A(n9031), .B(n3030), .Z(n7086) );
  HS65_LH_NAND2X4 U7699 ( .A(n6014), .B(n6013), .Z(n6018) );
  HS65_LH_NAND2X4 U7700 ( .A(n5903), .B(n5902), .Z(n5905) );
  HS65_LL_MUXI21X2 U7701 ( .D0(n3016), .D1(n3015), .S0(n3404), .Z(n4175) );
  HS65_LH_NOR2AX3 U7702 ( .A(n3024), .B(n3404), .Z(n3025) );
  HS65_LL_AND2X4 U7703 ( .A(n2962), .B(n2960), .Z(n2935) );
  HS65_LH_IVX4 U7704 ( .A(n6022), .Z(n6081) );
  HS65_LH_NAND2X4 U7705 ( .A(n5806), .B(n5805), .Z(n5810) );
  HS65_LL_AND2X4 U7706 ( .A(\u_DataPath/cw_memwb_i [2]), .B(n2960), .Z(n2961)
         );
  HS65_LH_MUXI21X5 U7707 ( .D0(n3098), .D1(n9377), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8427) );
  HS65_LL_NAND2X5 U7708 ( .A(n3030), .B(n2942), .Z(n7619) );
  HS65_LH_MUXI21X2 U7709 ( .D0(n3166), .D1(n9380), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8350) );
  HS65_LH_MUXI21X2 U7711 ( .D0(n8914), .D1(
        \u_DataPath/from_mem_data_out_i [28]), .S0(n3404), .Z(n8383) );
  HS65_LH_OAI12X3 U7713 ( .A(n5877), .B(n5874), .C(n5876), .Z(n5780) );
  HS65_LH_OAI12X3 U7714 ( .A(n6082), .B(n6019), .C(n6021), .Z(n6010) );
  HS65_LHS_XNOR2X3 U7715 ( .A(n8687), .B(n3126), .Z(\u_DataPath/pc_4_i [3]) );
  HS65_LH_OAI12X3 U7716 ( .A(n5871), .B(n5775), .C(n5777), .Z(n5725) );
  HS65_LH_NOR2X3 U7718 ( .A(n7613), .B(n8932), .Z(n7616) );
  HS65_LH_BFX9 U7719 ( .A(n8286), .Z(n7890) );
  HS65_LH_OAI12X3 U7720 ( .A(n5897), .B(n5894), .C(n5896), .Z(n5719) );
  HS65_LH_BFX9 U7721 ( .A(n8283), .Z(n7883) );
  HS65_LH_NOR2X3 U7722 ( .A(n8163), .B(rst), .Z(\u_DataPath/rs_ex_i [0]) );
  HS65_LH_NOR2X3 U7723 ( .A(n2881), .B(rst), .Z(\u_DataPath/idex_rt_i [4]) );
  HS65_LH_OAI12X3 U7724 ( .A(n5891), .B(n5836), .C(n5838), .Z(n5833) );
  HS65_LH_NOR2X3 U7725 ( .A(n8184), .B(rst), .Z(\u_DataPath/idex_rt_i [2]) );
  HS65_LH_NOR2X3 U7726 ( .A(n8153), .B(rst), .Z(\u_DataPath/idex_rt_i [1]) );
  HS65_LH_OAI12X3 U7728 ( .A(n6100), .B(n6097), .C(n6099), .Z(n5921) );
  HS65_LH_OAI12X3 U7729 ( .A(n6094), .B(n6038), .C(n6040), .Z(n6035) );
  HS65_LH_OAI12X3 U7730 ( .A(n5885), .B(n5882), .C(n5884), .Z(n5721) );
  HS65_LH_IVX9 U7731 ( .A(n3470), .Z(n3416) );
  HS65_LH_OAI12X3 U7732 ( .A(n5863), .B(n5753), .C(n5755), .Z(n5727) );
  HS65_LL_OR2X4 U7733 ( .A(\u_DataPath/jaddr_i [19]), .B(n2881), .Z(n2880) );
  HS65_LH_NAND2X7 U7735 ( .A(n2983), .B(n2984), .Z(n7638) );
  HS65_LH_NAND2X4 U7736 ( .A(n5812), .B(n5811), .Z(n5816) );
  HS65_LL_NAND2AX4 U7737 ( .A(\u_DataPath/jaddr_i [20]), .B(n6339), .Z(n6332)
         );
  HS65_LH_BFX9 U7738 ( .A(n8283), .Z(n7884) );
  HS65_LH_NAND2AX7 U7739 ( .A(n8480), .B(n9151), .Z(n8263) );
  HS65_LH_NAND2AX7 U7740 ( .A(n8480), .B(n8910), .Z(n8231) );
  HS65_LH_OR2X9 U7741 ( .A(n9343), .B(n9217), .Z(n5805) );
  HS65_LH_NOR2X3 U7742 ( .A(n9235), .B(n8915), .Z(n2973) );
  HS65_LH_IVX9 U7744 ( .A(\u_DataPath/dataOut_exe_i [3]), .Z(n3307) );
  HS65_LHS_XNOR2X6 U7747 ( .A(\u_DataPath/jaddr_i [19]), .B(n9077), .Z(n7100)
         );
  HS65_LH_CNIVX3 U7748 ( .A(\u_DataPath/dataOut_exe_i [0]), .Z(n8131) );
  HS65_LL_IVX4 U7750 ( .A(\u_DataPath/cw_to_ex_i [3]), .Z(n5491) );
  HS65_LH_IVX4 U7752 ( .A(n9225), .Z(n7788) );
  HS65_LH_CNIVX3 U7753 ( .A(\u_DataPath/cw_to_ex_i [4]), .Z(n3448) );
  HS65_LH_OR2X9 U7754 ( .A(n9341), .B(n9220), .Z(n5811) );
  HS65_LL_IVX4 U7755 ( .A(\u_DataPath/cw_to_ex_i [2]), .Z(n5492) );
  HS65_LH_NOR2X5 U7757 ( .A(n9033), .B(n9215), .Z(n6097) );
  HS65_LH_NOR2X5 U7758 ( .A(n9039), .B(n9116), .Z(n6102) );
  HS65_LH_OR2X9 U7759 ( .A(n9341), .B(n9204), .Z(n5858) );
  HS65_LH_OR2X4 U7761 ( .A(n9035), .B(n9115), .Z(n5717) );
  HS65_LH_IVX9 U7762 ( .A(\u_DataPath/jaddr_i [18]), .Z(n8184) );
  HS65_LH_NOR2X5 U7765 ( .A(n8967), .B(n9220), .Z(n6066) );
  HS65_LH_NOR2X3 U7766 ( .A(n9077), .B(n9218), .Z(n6061) );
  HS65_LH_IVX9 U7767 ( .A(n8961), .Z(\u_DataPath/cw_memwb_i [2]) );
  HS65_LH_OR2X9 U7768 ( .A(n9342), .B(n9208), .Z(n5914) );
  HS65_LH_NOR2X5 U7769 ( .A(n9181), .B(n9226), .Z(n5960) );
  HS65_LH_IVX7 U7770 ( .A(n8682), .Z(n7667) );
  HS65_LH_IVX9 U7772 ( .A(n8700), .Z(n3120) );
  HS65_LLS_XNOR2X3 U7773 ( .A(n8966), .B(n8766), .Z(n2962) );
  HS65_LH_NOR2X5 U7774 ( .A(n9183), .B(n9232), .Z(n5976) );
  HS65_LH_NOR2X5 U7775 ( .A(n9171), .B(n9214), .Z(n5979) );
  HS65_LH_NOR2X5 U7777 ( .A(n9185), .B(n9230), .Z(n5990) );
  HS65_LH_IVX4 U7778 ( .A(n9222), .Z(n7715) );
  HS65_LL_NOR2AX3 U7781 ( .A(n3267), .B(n3814), .Z(n4919) );
  HS65_LL_NAND4ABX3 U7782 ( .A(n4603), .B(n4602), .C(n4601), .D(n4600), .Z(
        n4604) );
  HS65_LL_AO12X4 U7783 ( .A(n3030), .B(n8139), .C(n2947), .Z(n2948) );
  HS65_LLS_XNOR2X3 U7785 ( .A(n4248), .B(n4247), .Z(n4249) );
  HS65_LH_NOR2X2 U7786 ( .A(n9077), .B(n9218), .Z(n2875) );
  HS65_LH_CBI4I6X2 U7787 ( .A(n9346), .B(n5417), .C(n3529), .D(n2860), .Z(
        n3709) );
  HS65_LH_CNIVX3 U7788 ( .A(n9215), .Z(n7706) );
  HS65_LL_NOR2AX3 U7789 ( .A(n3472), .B(n3560), .Z(n5257) );
  HS65_LLS_XNOR2X3 U7790 ( .A(n8943), .B(n2847), .Z(n3053) );
  HS65_LLS_XNOR2X3 U7791 ( .A(n8151), .B(n7619), .Z(n7078) );
  HS65_LLS_XNOR2X3 U7792 ( .A(n8763), .B(n8969), .Z(n3035) );
  HS65_LL_AOI12X2 U7794 ( .A(n5297), .B(n5466), .C(n5300), .Z(n4685) );
  HS65_LL_NOR2X2 U7795 ( .A(n5041), .B(n4583), .Z(n3764) );
  HS65_LL_NAND3X2 U7796 ( .A(n5534), .B(n5533), .C(n5532), .Z(n5535) );
  HS65_LL_AOI12X2 U7797 ( .A(n4431), .B(n4204), .C(n4203), .Z(n4228) );
  HS65_LL_AND3X4 U7798 ( .A(n4708), .B(n5432), .C(n5416), .Z(n2904) );
  HS65_LLS_XNOR2X3 U7799 ( .A(n4021), .B(n4020), .Z(n5284) );
  HS65_LL_NAND2X2 U7800 ( .A(n3426), .B(n4839), .Z(n4432) );
  HS65_LL_OA22X4 U7801 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [30]), .C(
        n8380), .D(n3409), .Z(n2916) );
  HS65_LLS_XNOR2X3 U7802 ( .A(n4907), .B(n4906), .Z(n4908) );
  HS65_LLS_XNOR2X3 U7803 ( .A(n5613), .B(n5612), .Z(n5642) );
  HS65_LL_NOR2X2 U7804 ( .A(n4333), .B(n4328), .Z(n4304) );
  HS65_LL_NOR2AX3 U7805 ( .A(n4297), .B(n4296), .Z(n4298) );
  HS65_LL_NAND2X7 U7806 ( .A(n3230), .B(n3229), .Z(n5053) );
  HS65_LL_NAND3X2 U7807 ( .A(n5450), .B(n4996), .C(n5449), .Z(n4992) );
  HS65_LL_NOR2X3 U7808 ( .A(\lte_x_59/B[9] ), .B(n2871), .Z(n5396) );
  HS65_LH_CNIVX3 U7810 ( .A(n9231), .Z(n7783) );
  HS65_LL_NAND3X2 U7811 ( .A(n5534), .B(n5533), .C(n4988), .Z(n4989) );
  HS65_LL_IVX2 U7812 ( .A(n5355), .Z(n5467) );
  HS65_LL_AOI12X2 U7813 ( .A(n5068), .B(n5067), .C(n5066), .Z(n5069) );
  HS65_LH_AOI21X2 U7815 ( .A(\lte_x_59/B[28] ), .B(n4488), .C(n3447), .Z(n3453) );
  HS65_LH_CNIVX3 U7817 ( .A(n5081), .Z(n4990) );
  HS65_LH_OAI21X2 U7818 ( .A(n3515), .B(n4987), .C(n5529), .Z(n4988) );
  HS65_LH_CBI4I1X3 U7820 ( .A(n5587), .B(n5586), .C(n5585), .D(n5584), .Z(
        n5588) );
  HS65_LH_CBI4I1X3 U7821 ( .A(n5370), .B(n5369), .C(n5484), .D(n5368), .Z(
        n5371) );
  HS65_LH_CNIVX3 U7822 ( .A(n5482), .Z(n5353) );
  HS65_LHS_XOR2X3 U7823 ( .A(n4985), .B(\lte_x_59/B[16] ), .Z(n4857) );
  HS65_LH_NOR2X6 U7824 ( .A(n2840), .B(n5089), .Z(n3969) );
  HS65_LH_CNIVX3 U7825 ( .A(n3803), .Z(n3686) );
  HS65_LH_OAI21X3 U7826 ( .A(n4502), .B(n4889), .C(n4080), .Z(n4363) );
  HS65_LH_BFX9 U7827 ( .A(n6690), .Z(n7604) );
  HS65_LH_AOI22X1 U7828 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][27] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ), .D(
        n6362), .Z(n6208) );
  HS65_LH_AOI22X1 U7829 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][11] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ), .D(
        n6362), .Z(n6248) );
  HS65_LH_AOI22X1 U7831 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ), .B(n7525), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][26] ), .Z(n7325)
         );
  HS65_LH_AOI22X1 U7832 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][23] ), .D(
        n6362), .Z(n6228) );
  HS65_LH_AOI22X1 U7833 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][25] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ), .D(
        n6362), .Z(n7146) );
  HS65_LH_AOI22X1 U7834 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][28] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][28] ), .D(
        n7296), .Z(n6919) );
  HS65_LH_BFX9 U7835 ( .A(n6684), .Z(n7594) );
  HS65_LH_NOR2X6 U7836 ( .A(n6153), .B(n6152), .Z(n7296) );
  HS65_LH_AOI22X1 U7837 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][17] ), .B(n7525), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ), .Z(n6815)
         );
  HS65_LH_AOI22X1 U7838 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][17] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ), .D(
        n2891), .Z(n6810) );
  HS65_LH_AOI22X1 U7839 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][18] ), .D(
        n7296), .Z(n6662) );
  HS65_LH_BFX9 U7840 ( .A(n6753), .Z(n7524) );
  HS65_LH_AOI22X1 U7841 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ), .B(n7525), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ), .Z(n6835)
         );
  HS65_LH_AO22X4 U7842 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ), .D(n7318), .Z(n6832) );
  HS65_LH_BFX9 U7843 ( .A(n7295), .Z(n6941) );
  HS65_LH_AOI22X1 U7844 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][31] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ), .D(
        n7296), .Z(n6879) );
  HS65_LH_NOR2X6 U7845 ( .A(n6348), .B(n6333), .Z(n7320) );
  HS65_LL_NOR2AX3 U7847 ( .A(n3075), .B(n3074), .Z(n3077) );
  HS65_LH_AOI312X2 U7848 ( .A(opcode_i[1]), .B(n7777), .C(n7693), .D(n9082), 
        .E(n7692), .F(n7691), .Z(n8102) );
  HS65_LH_OAI21X2 U7849 ( .A(n7697), .B(n8055), .C(n9082), .Z(n7683) );
  HS65_LH_CNIVX3 U7850 ( .A(n4655), .Z(n4656) );
  HS65_LH_CBI4I6X2 U7851 ( .A(n5549), .B(n5548), .C(n5547), .D(n5546), .Z(
        n5553) );
  HS65_LL_NOR2AX3 U7852 ( .A(n5504), .B(n5571), .Z(n5574) );
  HS65_LL_NOR2AX3 U7853 ( .A(n2853), .B(n5567), .Z(n5343) );
  HS65_LH_NOR2X2 U7854 ( .A(n4973), .B(n4972), .Z(n4975) );
  HS65_LH_AOI22X1 U7855 ( .A(n4717), .B(n4715), .C(n4714), .D(n3133), .Z(n4716) );
  HS65_LH_CBI4I6X2 U7856 ( .A(n5332), .B(n5331), .C(n5330), .D(n5329), .Z(
        n5337) );
  HS65_LH_NAND3X2 U7857 ( .A(n5328), .B(n5327), .C(n5326), .Z(n5329) );
  HS65_LH_NAND2X2 U7858 ( .A(n9376), .B(n8549), .Z(n3162) );
  HS65_LL_NAND2AX4 U7859 ( .A(n3588), .B(n3587), .Z(n3589) );
  HS65_LH_OAI22X1 U7860 ( .A(n5041), .B(n4583), .C(n3756), .D(n4796), .Z(n4463) );
  HS65_LH_NOR2AX3 U7861 ( .A(n2864), .B(n5004), .Z(n3841) );
  HS65_LH_NOR2X2 U7862 ( .A(n9346), .B(n4724), .Z(n3424) );
  HS65_LH_NOR4ABX2 U7863 ( .A(n5293), .B(n5275), .C(n5360), .D(n5354), .Z(
        n5341) );
  HS65_LH_CNIVX3 U7864 ( .A(n5352), .Z(n5288) );
  HS65_LHS_XOR2X3 U7865 ( .A(\lte_x_59/B[7] ), .B(n5030), .Z(n4771) );
  HS65_LH_CNIVX3 U7866 ( .A(n4876), .Z(n4877) );
  HS65_LL_NAND4ABX3 U7867 ( .A(n3841), .B(n3840), .C(n3839), .D(n3838), .Z(
        n4835) );
  HS65_LH_NAND2X7 U7869 ( .A(n7665), .B(n7646), .Z(n7653) );
  HS65_LH_CNIVX3 U7870 ( .A(n3629), .Z(n3630) );
  HS65_LH_AOI22X1 U7872 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ), .B(n7604), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ), .Z(n7464)
         );
  HS65_LH_AOI22X1 U7873 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ), .D(
        n6362), .Z(n6308) );
  HS65_LH_AOI22X1 U7874 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ), .Z(n7376)
         );
  HS65_LH_AOI22X1 U7875 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ), .B(n7525), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][3] ), .Z(n7395)
         );
  HS65_LH_AOI22X1 U7876 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][10] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][10] ), .Z(n7213)
         );
  HS65_LH_AO22X4 U7877 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ), .B(n2891), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ), .D(
        n7415), .Z(n7418) );
  HS65_LH_AOI22X1 U7878 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][13] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ), .D(
        n6362), .Z(n7164) );
  HS65_LH_AOI22X1 U7879 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ), .B(n7604), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ), .Z(n7530)
         );
  HS65_LH_CBI4I1X3 U7880 ( .A(n5648), .B(n5422), .C(n4488), .D(
        \sub_x_53/A[29] ), .Z(n4361) );
  HS65_LH_AOI22X1 U7882 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ), .D(
        n6362), .Z(n6188) );
  HS65_LH_AOI22X1 U7883 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ), .B(n7604), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][21] ), .Z(n7605)
         );
  HS65_LH_AOI22X1 U7884 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ), .Z(n7595)
         );
  HS65_LH_AOI22X1 U7885 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ), .Z(n6708)
         );
  HS65_LH_AOI22X1 U7886 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][24] ), .D(
        n6362), .Z(n6288) );
  HS65_LH_AOI22X1 U7887 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ), .B(n7604), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ), .Z(n7570)
         );
  HS65_LH_AOI22X1 U7888 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][28] ), .B(n7525), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ), .Z(n7500)
         );
  HS65_LH_AOI22X1 U7889 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ), .B(n7604), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][28] ), .Z(n7504)
         );
  HS65_LH_AOI22X1 U7890 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ), .B(n7604), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ), .Z(n7550)
         );
  HS65_LH_AOI22X1 U7891 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ), .Z(n7546)
         );
  HS65_LH_AOI22X1 U7892 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][6] ), .Z(n7253)
         );
  HS65_LH_BFX9 U7893 ( .A(n7319), .Z(n7586) );
  HS65_LH_BFX9 U7894 ( .A(n7329), .Z(n7599) );
  HS65_LH_BFX9 U7895 ( .A(n7331), .Z(n7601) );
  HS65_LH_AOI22X1 U7896 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ), .B(n7604), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ), .Z(n7444)
         );
  HS65_LH_AOI22X1 U7897 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][0] ), .Z(n7441)
         );
  HS65_LH_NOR2X2 U7898 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .B(n8157), 
        .Z(n8122) );
  HS65_LH_NAND2X2 U7899 ( .A(\u_DataPath/jaddr_i [22]), .B(n8163), .Z(n6146)
         );
  HS65_LH_AO22X4 U7905 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ), .D(
        n7292), .Z(n6219) );
  HS65_LH_AOI22X1 U7906 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][27] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ), .D(
        n7296), .Z(n6217) );
  HS65_LH_AO22X4 U7907 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][27] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][27] ), .D(
        n6382), .Z(n6220) );
  HS65_LH_AO22X4 U7908 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ), .D(
        n6635), .Z(n6216) );
  HS65_LH_AOI22X1 U7909 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ), .D(
        n6172), .Z(n6213) );
  HS65_LH_AO22X4 U7910 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][27] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ), .D(
        n6619), .Z(n6205) );
  HS65_LH_AOI22X1 U7911 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ), .D(
        n6363), .Z(n6207) );
  HS65_LH_AO22X4 U7912 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][27] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][27] ), .D(
        n6629), .Z(n6209) );
  HS65_LH_AO22X4 U7913 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][27] ), .D(
        n6627), .Z(n6210) );
  HS65_LH_AOI22X1 U7914 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][15] ), .D(
        n2888), .Z(n6368) );
  HS65_LH_AOI22X1 U7915 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][15] ), .D(
        n7272), .Z(n6374) );
  HS65_LH_AOI22X1 U7916 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][15] ), .D(
        n6600), .Z(n6375) );
  HS65_LH_AO22X4 U7917 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][15] ), .D(
        n7276), .Z(n6372) );
  HS65_LH_AO22X4 U7918 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][15] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][15] ), .D(
        n6383), .Z(n6388) );
  HS65_LH_AO22X4 U7919 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ), .D(
        n7284), .Z(n6380) );
  HS65_LH_AOI22X1 U7920 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ), .D(
        n7296), .Z(n6257) );
  HS65_LH_AO22X4 U7921 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][11] ), .D(
        n6382), .Z(n6260) );
  HS65_LH_AO22X4 U7922 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ), .D(
        n6635), .Z(n6256) );
  HS65_LH_AOI22X1 U7923 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][11] ), .D(
        n6172), .Z(n6253) );
  HS65_LH_AO22X4 U7924 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][11] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ), .D(
        n6619), .Z(n6245) );
  HS65_LH_AO22X4 U7925 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][11] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][11] ), .D(
        n6629), .Z(n6249) );
  HS65_LH_AO22X4 U7926 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][11] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ), .D(
        n6627), .Z(n6250) );
  HS65_LH_AOI22X1 U7927 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ), .D(
        n2888), .Z(n6517) );
  HS65_LH_AOI22X1 U7928 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][19] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][19] ), .D(
        n7272), .Z(n6521) );
  HS65_LH_AOI22X1 U7929 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][19] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][19] ), .D(
        n6600), .Z(n6522) );
  HS65_LH_AO22X4 U7930 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][19] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][19] ), .D(
        n7276), .Z(n6519) );
  HS65_LH_AO22X4 U7931 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][19] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ), .D(
        n6383), .Z(n6529) );
  HS65_LH_AOI22X1 U7932 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][19] ), .D(
        n6171), .Z(n6524) );
  HS65_LH_AO22X4 U7933 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ), .D(
        n7284), .Z(n6525) );
  HS65_LH_AOI22X1 U7934 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][3] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][3] ), .D(
        n2888), .Z(n6577) );
  HS65_LH_AOI22X1 U7935 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][3] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ), .D(
        n6625), .Z(n6581) );
  HS65_LH_AOI22X1 U7936 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ), .D(
        n6600), .Z(n6582) );
  HS65_LH_AO22X4 U7937 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][3] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ), .D(
        n7276), .Z(n6579) );
  HS65_LH_AO22X4 U7938 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ), .D(
        n6383), .Z(n6589) );
  HS65_LH_AOI22X1 U7939 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][3] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ), .D(
        n6171), .Z(n6584) );
  HS65_LH_AO22X4 U7940 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][3] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ), .D(
        n7282), .Z(n6586) );
  HS65_LH_AOI22X1 U7941 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ), .D(
        n2888), .Z(n6396) );
  HS65_LH_AOI22X1 U7942 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ), .D(
        n7272), .Z(n6400) );
  HS65_LH_AOI22X1 U7943 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ), .D(
        n6600), .Z(n6401) );
  HS65_LH_AO22X4 U7944 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ), .D(
        n7276), .Z(n6398) );
  HS65_LH_AO22X4 U7945 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][10] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][10] ), .D(
        n6383), .Z(n6408) );
  HS65_LH_AO22X4 U7946 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ), .D(
        n7284), .Z(n6404) );
  HS65_LH_AOI22X1 U7947 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ), .D(
        n2888), .Z(n6497) );
  HS65_LH_AOI22X1 U7948 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][26] ), .D(
        n7272), .Z(n6501) );
  HS65_LH_AOI22X1 U7949 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][26] ), .D(
        n6600), .Z(n6502) );
  HS65_LH_AO22X4 U7950 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][26] ), .D(
        n7276), .Z(n6499) );
  HS65_LH_AO22X4 U7951 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][26] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ), .D(
        n6383), .Z(n6509) );
  HS65_LH_AOI22X1 U7952 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][26] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ), .D(
        n6171), .Z(n6504) );
  HS65_LH_AO22X4 U7953 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ), .D(
        n7284), .Z(n6505) );
  HS65_LH_AOI22X1 U7954 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][26] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ), .D(n6746), 
        .Z(n7324) );
  HS65_LH_AO22X4 U7955 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ), .D(
        n7319), .Z(n7321) );
  HS65_LH_AOI22X1 U7956 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ), .D(
        n6670), .Z(n7316) );
  HS65_LH_AOI22X1 U7957 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][26] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][26] ), .D(n6740), 
        .Z(n7315) );
  HS65_LH_AO22X4 U7958 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][26] ), .B(n7578), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ), .Z(n7314)
         );
  HS65_LH_AO22X4 U7959 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ), .B(n9373), 
        .C(n7311), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ), .Z(n7313)
         );
  HS65_LH_AO22X4 U7960 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][26] ), .B(n7523), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][26] ), .Z(n7327)
         );
  HS65_LH_AOI22X1 U7961 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][26] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ), .Z(n7326)
         );
  HS65_LH_AO22X4 U7962 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][26] ), .Z(n7337)
         );
  HS65_LH_AO22X4 U7963 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][26] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][26] ), .Z(n7338)
         );
  HS65_LH_AOI22X1 U7964 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ), .D(
        n7296), .Z(n6237) );
  HS65_LH_AO22X4 U7965 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ), .D(
        n6382), .Z(n6240) );
  HS65_LH_AO22X4 U7966 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][23] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ), .D(
        n6635), .Z(n6236) );
  HS65_LH_AOI22X1 U7967 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ), .D(
        n6172), .Z(n6233) );
  HS65_LH_AO22X4 U7968 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][23] ), .D(
        n6619), .Z(n6225) );
  HS65_LH_AO22X4 U7969 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ), .D(
        n6629), .Z(n6229) );
  HS65_LH_AO22X4 U7970 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ), .D(
        n6627), .Z(n6230) );
  HS65_LH_AOI22X1 U7971 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ), .D(
        n2888), .Z(n6537) );
  HS65_LH_AOI22X1 U7972 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][12] ), .D(
        n6625), .Z(n6541) );
  HS65_LH_AOI22X1 U7973 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][12] ), .D(
        n6600), .Z(n6542) );
  HS65_LH_AO22X4 U7974 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][12] ), .D(
        n7276), .Z(n6539) );
  HS65_LH_AO22X4 U7975 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][12] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][12] ), .D(
        n6383), .Z(n6549) );
  HS65_LH_AOI22X1 U7976 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][12] ), .D(
        n6171), .Z(n6544) );
  HS65_LH_AO22X4 U7977 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ), .D(
        n7284), .Z(n6545) );
  HS65_LH_AOI22X1 U7978 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ), .D(
        n2888), .Z(n6437) );
  HS65_LH_AOI22X1 U7979 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ), .D(
        n7272), .Z(n6441) );
  HS65_LH_AOI22X1 U7980 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ), .D(
        n6600), .Z(n6442) );
  HS65_LH_AO22X4 U7981 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ), .D(
        n7276), .Z(n6439) );
  HS65_LH_AO22X4 U7982 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][7] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ), .D(
        n6383), .Z(n6449) );
  HS65_LH_AOI22X1 U7983 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ), .D(
        n6171), .Z(n6444) );
  HS65_LH_AO22X4 U7984 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][7] ), .D(
        n7284), .Z(n6445) );
  HS65_LH_AOI22X1 U7985 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][29] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][29] ), .D(
        n7272), .Z(n7280) );
  HS65_LH_AOI22X1 U7986 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][29] ), .D(
        n6600), .Z(n7281) );
  HS65_LH_AO22X4 U7987 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ), .D(
        n7284), .Z(n7289) );
  HS65_LH_AOI22X1 U7988 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ), .D(
        n6172), .Z(n7287) );
  HS65_LH_AO22X4 U7989 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][29] ), .D(
        n7292), .Z(n7300) );
  HS65_LH_AOI22X1 U7990 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][29] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ), .D(
        n7296), .Z(n7298) );
  HS65_LH_AOI22X1 U7991 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ), .D(
        n7272), .Z(n6935) );
  HS65_LH_AOI22X1 U7992 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ), .D(
        n6600), .Z(n6936) );
  HS65_LH_AO22X4 U7993 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][5] ), .D(
        n7284), .Z(n6939) );
  HS65_LH_AOI22X1 U7994 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ), .D(
        n6172), .Z(n6937) );
  HS65_LH_AO22X4 U7995 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][5] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ), .D(n6382), .Z(n6946) );
  HS65_LH_AO22X4 U7996 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][5] ), .D(
        n6383), .Z(n6945) );
  HS65_LH_AO22X4 U7997 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][25] ), .D(
        n7171), .Z(n2883) );
  HS65_LH_AO22X4 U7998 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ), .D(
        n6635), .Z(n7152) );
  HS65_LH_AO22X4 U7999 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ), .D(
        n6637), .Z(n7151) );
  HS65_LH_AO22X4 U8000 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][25] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ), .D(
        n7285), .Z(n2882) );
  HS65_LH_AO22X4 U8001 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][25] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ), .D(
        n6627), .Z(n7148) );
  HS65_LH_AOI22X1 U8002 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ), .D(
        n7296), .Z(n7153) );
  HS65_LH_AO22X4 U8003 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][25] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ), .D(
        n6619), .Z(n7143) );
  HS65_LH_AOI22X1 U8004 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][9] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ), .D(
        n6362), .Z(n7126) );
  HS65_LH_AO22X4 U8005 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ), .D(n6619), .Z(n7123) );
  HS65_LH_AO22X4 U8006 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][9] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ), .D(
        n6627), .Z(n7128) );
  HS65_LH_AO22X4 U8007 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ), .D(
        n6635), .Z(n7134) );
  HS65_LH_AOI22X1 U8008 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ), .D(n7296), .Z(n7135) );
  HS65_LH_AOI22X1 U8009 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][28] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ), .D(
        n6624), .Z(n6914) );
  HS65_LH_AO22X4 U8010 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ), .D(
        n7284), .Z(n6917) );
  HS65_LH_AOI22X1 U8011 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][28] ), .D(
        n6172), .Z(n6915) );
  HS65_LH_AOI22X1 U8012 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][4] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ), .D(
        n7272), .Z(n6632) );
  HS65_LH_AOI22X1 U8013 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][4] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ), .D(
        n6600), .Z(n6633) );
  HS65_LH_AO22X4 U8014 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ), .D(
        n7284), .Z(n6640) );
  HS65_LH_AOI22X1 U8015 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ), .D(
        n6172), .Z(n6638) );
  HS65_LH_AOI22X1 U8016 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ), .D(n7296), .Z(n6642) );
  HS65_LH_AO22X4 U8017 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ), .D(
        n7292), .Z(n6644) );
  HS65_LH_AOI22X1 U8018 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][4] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ), .D(
        n6362), .Z(n6623) );
  HS65_LH_AOI22X1 U8019 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ), .D(
        n2888), .Z(n6457) );
  HS65_LH_AOI22X1 U8020 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][8] ), .D(
        n7272), .Z(n6461) );
  HS65_LH_AO22X4 U8021 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][8] ), .D(
        n7276), .Z(n6459) );
  HS65_LH_AO22X4 U8022 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][8] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ), .D(
        n6383), .Z(n6469) );
  HS65_LH_AOI22X1 U8023 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ), .D(
        n6171), .Z(n6464) );
  HS65_LH_AO22X4 U8024 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][8] ), .D(
        n7284), .Z(n6465) );
  HS65_LH_AOI22X1 U8025 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][20] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ), .D(
        n6624), .Z(n6854) );
  HS65_LH_AO22X4 U8026 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ), .D(
        n7284), .Z(n6857) );
  HS65_LH_AOI22X1 U8027 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ), .D(
        n6172), .Z(n6855) );
  HS65_LH_AOI22X1 U8028 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][16] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ), .D(
        n7296), .Z(n6177) );
  HS65_LH_AO22X4 U8029 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][16] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][16] ), .D(
        n6382), .Z(n6180) );
  HS65_LH_AO22X4 U8030 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ), .D(
        n6635), .Z(n6176) );
  HS65_LH_AOI22X1 U8031 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][16] ), .D(
        n6172), .Z(n6173) );
  HS65_LH_AOI22X1 U8032 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][16] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ), .D(
        n6171), .Z(n6174) );
  HS65_LH_AO22X4 U8033 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][16] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ), .D(
        n6619), .Z(n6163) );
  HS65_LH_AOI22X1 U8034 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ), .D(
        n6363), .Z(n6165) );
  HS65_LH_AO22X4 U8035 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][16] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][16] ), .D(
        n6629), .Z(n6167) );
  HS65_LH_AO22X4 U8036 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][16] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][16] ), .D(
        n6627), .Z(n6168) );
  HS65_LH_AOI22X1 U8037 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ), .D(
        n7272), .Z(n6893) );
  HS65_LH_AO22X4 U8038 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ), .D(
        n7284), .Z(n6897) );
  HS65_LH_AOI22X1 U8039 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][17] ), .D(
        n6172), .Z(n6895) );
  HS65_LH_AO22X4 U8040 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][17] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ), .D(
        n6382), .Z(n6902) );
  HS65_LH_AO22X4 U8041 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][17] ), .D(
        n6383), .Z(n6901) );
  HS65_LH_AO22X4 U8042 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][17] ), .D(
        n7318), .Z(n6812) );
  HS65_LH_AO22X4 U8043 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][17] ), .D(
        n7319), .Z(n6811) );
  HS65_LH_AOI22X1 U8044 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ), .Z(n6820)
         );
  HS65_LH_AOI22X1 U8045 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ), .Z(n6819)
         );
  HS65_LH_AO22X4 U8046 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ), .Z(n6822)
         );
  HS65_LH_AO22X4 U8047 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ), .Z(n6821)
         );
  HS65_LH_AO22X4 U8048 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][17] ), .B(n7523), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][17] ), .Z(n6817)
         );
  HS65_LH_AOI22X1 U8049 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][17] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][17] ), .Z(n6816)
         );
  HS65_LH_AO22X4 U8050 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ), .B(n9373), 
        .C(n7311), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][17] ), .Z(n6807)
         );
  HS65_LH_AO22X4 U8051 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][17] ), .B(n7429), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ), .Z(n6808)
         );
  HS65_LH_AOI22X1 U8052 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][17] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][17] ), .D(n6740), 
        .Z(n6809) );
  HS65_LH_AOI22X1 U8053 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ), .D(
        n2888), .Z(n6557) );
  HS65_LH_AOI22X1 U8054 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][2] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ), .D(
        n7272), .Z(n6561) );
  HS65_LH_AO22X4 U8055 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ), .D(
        n6383), .Z(n6569) );
  HS65_LH_AO22X4 U8056 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ), .D(
        n6637), .Z(n6565) );
  HS65_LH_AOI22X1 U8057 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][18] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][18] ), .D(
        n7272), .Z(n6656) );
  HS65_LH_AOI22X1 U8058 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][18] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][18] ), .D(
        n6624), .Z(n6657) );
  HS65_LH_AO22X4 U8059 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ), .D(
        n7284), .Z(n6660) );
  HS65_LH_AOI22X1 U8060 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][18] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ), .D(
        n6362), .Z(n6653) );
  HS65_LH_AO22X4 U8061 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ), .D(
        n6382), .Z(n6665) );
  HS65_LH_AO22X4 U8062 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][18] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][18] ), .D(
        n6383), .Z(n6664) );
  HS65_LH_AOI22X1 U8063 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ), .D(
        n2888), .Z(n6598) );
  HS65_LH_AOI22X1 U8064 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ), .D(
        n6625), .Z(n6603) );
  HS65_LH_AO22X4 U8065 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ), .D(
        n6627), .Z(n6602) );
  HS65_LH_AO22X4 U8066 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][1] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][1] ), .D(
        n6383), .Z(n6611) );
  HS65_LH_AO22X4 U8067 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ), .D(
        n6637), .Z(n6607) );
  HS65_LH_AO22X4 U8068 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ), .D(
        n6635), .Z(n6608) );
  HS65_LH_AOI22X1 U8069 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][1] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ), .D(
        n6171), .Z(n6606) );
  HS65_LH_AOI22X1 U8070 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][1] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][1] ), .D(
        n6670), .Z(n6830) );
  HS65_LH_AOI22X1 U8071 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][1] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][1] ), .D(n6740), 
        .Z(n6829) );
  HS65_LH_AO22X4 U8072 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][1] ), .B(n7429), 
        .C(n6952), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][1] ), .Z(n6828) );
  HS65_LH_AO22X4 U8073 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ), .B(n9373), 
        .C(n7311), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ), .Z(n6827) );
  HS65_LH_AOI22X1 U8074 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][1] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ), .Z(n6840)
         );
  HS65_LH_AOI22X1 U8075 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][1] ), .Z(n6839)
         );
  HS65_LH_AO22X4 U8076 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][1] ), .Z(n6842)
         );
  HS65_LH_AO22X4 U8077 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][1] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ), .Z(n6841)
         );
  HS65_LH_AOI22X1 U8078 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][1] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][1] ), .Z(n6836)
         );
  HS65_LH_AO22X4 U8079 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][1] ), .D(
        n7319), .Z(n6831) );
  HS65_LH_AOI22X1 U8080 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][0] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ), .D(
        n2888), .Z(n6416) );
  HS65_LH_AOI22X1 U8081 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][0] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][0] ), .D(
        n7272), .Z(n6420) );
  HS65_LH_AO22X4 U8082 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][0] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][0] ), .D(
        n7276), .Z(n6418) );
  HS65_LH_AO22X4 U8083 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][0] ), .D(
        n6383), .Z(n6429) );
  HS65_LH_AOI22X1 U8084 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][0] ), .D(
        n6171), .Z(n6423) );
  HS65_LH_AO22X4 U8085 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ), .D(
        n7284), .Z(n6424) );
  HS65_LH_NOR2X2 U8086 ( .A(n7738), .B(n7775), .Z(n7763) );
  HS65_LH_CBI4I1X3 U8087 ( .A(n8098), .B(n8122), .C(n8097), .D(n8635), .Z(
        n8099) );
  HS65_LH_AO22X4 U8088 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][31] ), .D(
        n7284), .Z(n6877) );
  HS65_LH_AOI22X1 U8089 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ), .D(
        n6172), .Z(n6875) );
  HS65_LH_AO22X4 U8090 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][31] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ), .D(
        n6382), .Z(n6882) );
  HS65_LH_AO22X4 U8091 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][31] ), .D(
        n6383), .Z(n6881) );
  HS65_LH_NOR2X2 U8093 ( .A(n2842), .B(n5376), .Z(n5404) );
  HS65_LH_NAND2X2 U8094 ( .A(n5105), .B(n5104), .Z(n5052) );
  HS65_LH_OAI21X2 U8095 ( .A(n5313), .B(n5299), .C(n5055), .Z(n5058) );
  HS65_LH_NAND2X2 U8096 ( .A(n5054), .B(n5053), .Z(n5055) );
  HS65_LH_NAND2X2 U8097 ( .A(n4676), .B(n5061), .Z(n5065) );
  HS65_LH_NOR2X2 U8098 ( .A(n5062), .B(n3272), .Z(n5064) );
  HS65_LH_NOR2X2 U8099 ( .A(n5300), .B(n5047), .Z(n5056) );
  HS65_LH_NOR2X2 U8100 ( .A(n5105), .B(n5104), .Z(n5047) );
  HS65_LH_NOR2X2 U8101 ( .A(n5083), .B(n5064), .Z(n5067) );
  HS65_LH_NOR2X2 U8102 ( .A(n5004), .B(n5231), .Z(n5357) );
  HS65_LH_NOR2X2 U8103 ( .A(\lte_x_59/B[3] ), .B(n5089), .Z(n5383) );
  HS65_LH_NOR2X2 U8104 ( .A(n5136), .B(n4660), .Z(n5091) );
  HS65_LH_NOR2X2 U8105 ( .A(n5652), .B(n5654), .Z(n5361) );
  HS65_LH_NOR2X2 U8106 ( .A(n2849), .B(n3372), .Z(n5430) );
  HS65_LH_NAND2X2 U8107 ( .A(\lte_x_59/B[3] ), .B(n5089), .Z(n5090) );
  HS65_LH_NOR2X2 U8108 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n7834), .Z(n5570)
         );
  HS65_LH_CNIVX3 U8109 ( .A(n5564), .Z(n5565) );
  HS65_LH_CNIVX3 U8110 ( .A(n5325), .Z(n5326) );
  HS65_LH_NAND2X2 U8111 ( .A(n5041), .B(n5040), .Z(n5328) );
  HS65_LH_AOI21X2 U8112 ( .A(n5549), .B(n5547), .C(n5465), .Z(n5331) );
  HS65_LH_NOR2X2 U8113 ( .A(n4575), .B(n5383), .Z(n5385) );
  HS65_LH_OAI12X3 U8114 ( .A(n4817), .B(n5382), .C(n4819), .Z(n5386) );
  HS65_LH_NOR2X2 U8115 ( .A(n5123), .B(\sub_x_53/A[0] ), .Z(n5382) );
  HS65_LH_NOR2X2 U8116 ( .A(n5380), .B(n4637), .Z(n5390) );
  HS65_LH_NOR2X2 U8117 ( .A(n2865), .B(\lte_x_59/B[6] ), .Z(n5380) );
  HS65_LH_NOR2X2 U8118 ( .A(n5388), .B(n4100), .Z(n5381) );
  HS65_LH_NAND2X2 U8119 ( .A(\lte_x_59/B[8] ), .B(n3360), .Z(n5397) );
  HS65_LH_NAND2X2 U8120 ( .A(\lte_x_59/B[9] ), .B(n2871), .Z(n5395) );
  HS65_LH_OAI21X2 U8121 ( .A(n5405), .B(n5404), .C(n4050), .Z(n5409) );
  HS65_LH_OAI21X2 U8122 ( .A(n4915), .B(n5406), .C(n3893), .Z(n5407) );
  HS65_LH_OAI21X2 U8123 ( .A(n5400), .B(n5399), .C(n4013), .Z(n5401) );
  HS65_LH_NOR2X2 U8124 ( .A(n5404), .B(n5377), .Z(n5378) );
  HS65_LH_NOR2X2 U8125 ( .A(n3521), .B(n3365), .Z(n5377) );
  HS65_LH_OAI21X2 U8126 ( .A(n5272), .B(n5430), .C(n5270), .Z(n5431) );
  HS65_LH_OAI21X2 U8127 ( .A(n5506), .B(n3515), .C(n5531), .Z(n5433) );
  HS65_LH_OAI21X2 U8128 ( .A(n4418), .B(n4407), .C(n5434), .Z(n5438) );
  HS65_LH_NAND2X2 U8129 ( .A(\sub_x_53/A[29] ), .B(n5447), .Z(n5448) );
  HS65_LH_NAND2X2 U8130 ( .A(\sub_x_53/A[27] ), .B(n3385), .Z(n5443) );
  HS65_LH_NOR2X2 U8131 ( .A(n5419), .B(n4407), .Z(n5420) );
  HS65_LH_NOR2X2 U8132 ( .A(\sub_x_53/A[20] ), .B(n3376), .Z(n5419) );
  HS65_LH_NAND2X2 U8134 ( .A(n5514), .B(n4672), .Z(n5303) );
  HS65_LH_NAND2X2 U8135 ( .A(n5270), .B(n4244), .Z(n5533) );
  HS65_LH_NAND2X2 U8137 ( .A(n5022), .B(n5021), .Z(n5003) );
  HS65_LH_NAND2X2 U8138 ( .A(n4984), .B(n5001), .Z(n5002) );
  HS65_LH_OAI21X2 U8139 ( .A(n5357), .B(n5006), .C(n5534), .Z(n5007) );
  HS65_LH_NAND2X2 U8140 ( .A(n4986), .B(n5005), .Z(n5006) );
  HS65_LH_OAI21X2 U8141 ( .A(n5344), .B(n5347), .C(n5564), .Z(n5013) );
  HS65_LH_NOR2X2 U8142 ( .A(n5342), .B(n5503), .Z(n5015) );
  HS65_LH_OAI21X3 U8143 ( .A(n5192), .B(n5012), .C(n5289), .Z(n5580) );
  HS65_LH_AOI21X2 U8144 ( .A(n5098), .B(n5552), .C(n5043), .Z(n5044) );
  HS65_LH_OAI21X2 U8145 ( .A(n5327), .B(n5095), .C(n5544), .Z(n5043) );
  HS65_LH_NAND2X2 U8146 ( .A(n5552), .B(n5034), .Z(n5046) );
  HS65_LH_NOR2X2 U8147 ( .A(n5042), .B(n5033), .Z(n5034) );
  HS65_LH_AOI21X2 U8148 ( .A(n5039), .B(n5038), .C(n5554), .Z(n5045) );
  HS65_LH_NOR2X2 U8149 ( .A(n5036), .B(n5037), .Z(n5038) );
  HS65_LH_OAI21X2 U8150 ( .A(n5549), .B(n5548), .C(n5547), .Z(n5039) );
  HS65_LH_OAI21X2 U8151 ( .A(n5052), .B(n5300), .C(n5297), .Z(n5060) );
  HS65_LH_OAI21X2 U8153 ( .A(n5516), .B(n5514), .C(n5517), .Z(n5068) );
  HS65_LH_NAND2X2 U8154 ( .A(n5062), .B(n3272), .Z(n5063) );
  HS65_LH_NAND2X2 U8155 ( .A(n5540), .B(n5056), .Z(n5051) );
  HS65_LH_NAND2X2 U8156 ( .A(n5050), .B(n5067), .Z(n5071) );
  HS65_LH_NOR2X2 U8157 ( .A(n5049), .B(n5514), .Z(n5050) );
  HS65_LH_NOR2X2 U8158 ( .A(n4671), .B(n5048), .Z(n5049) );
  HS65_LH_NOR2X2 U8159 ( .A(n5022), .B(n5021), .Z(n5024) );
  HS65_LH_NOR2X2 U8160 ( .A(n4984), .B(n5001), .Z(n5023) );
  HS65_LH_NOR2X2 U8161 ( .A(n5357), .B(n5355), .Z(n5025) );
  HS65_LH_NAND3X2 U8163 ( .A(n5540), .B(n5405), .C(n4050), .Z(n5099) );
  HS65_LH_OAI21X2 U8164 ( .A(n5093), .B(n5092), .C(n5552), .Z(n5094) );
  HS65_LH_NOR2X2 U8165 ( .A(n5548), .B(n5091), .Z(n5093) );
  HS65_LH_NAND3X2 U8166 ( .A(n5318), .B(n5547), .C(n5317), .Z(n5092) );
  HS65_LH_NOR2X2 U8167 ( .A(n2860), .B(n4967), .Z(n4968) );
  HS65_LH_CNIVX3 U8168 ( .A(n5142), .Z(n5147) );
  HS65_LH_OAI21X2 U8170 ( .A(n5130), .B(n5129), .C(n5128), .Z(n5132) );
  HS65_LHS_XNOR2X3 U8171 ( .A(\lte_x_59/B[28] ), .B(n5423), .Z(n4761) );
  HS65_LH_NAND2X2 U8172 ( .A(\lte_x_59/B[7] ), .B(n4351), .Z(n3524) );
  HS65_LH_NOR2X2 U8173 ( .A(n4682), .B(n4583), .Z(n3525) );
  HS65_LH_AND2X4 U8174 ( .A(n9376), .B(n8499), .Z(n3322) );
  HS65_LH_AOI21X2 U8176 ( .A(n3446), .B(n3445), .C(n5646), .Z(n3447) );
  HS65_LH_CNIVX3 U8177 ( .A(n3834), .Z(n3446) );
  HS65_LH_NOR2X2 U8178 ( .A(n5373), .B(n4682), .Z(n5311) );
  HS65_LH_NAND2X2 U8180 ( .A(n2843), .B(n4683), .Z(n5297) );
  HS65_LH_NAND2X2 U8181 ( .A(\lte_x_59/B[7] ), .B(n5312), .Z(n4663) );
  HS65_LH_NAND2X2 U8182 ( .A(n2865), .B(\lte_x_59/B[6] ), .Z(n4664) );
  HS65_LH_CBI4I6X2 U8183 ( .A(n5387), .B(n5388), .C(n4143), .D(n4666), .Z(
        n4667) );
  HS65_LH_AND3X4 U8185 ( .A(n5322), .B(n4658), .C(n5317), .Z(n4659) );
  HS65_LH_CNIVX3 U8186 ( .A(n5388), .Z(n4658) );
  HS65_LH_CNIVX3 U8187 ( .A(n5583), .Z(n5587) );
  HS65_LH_CNIVX3 U8188 ( .A(n5544), .Z(n5558) );
  HS65_LH_CNIVX3 U8189 ( .A(n5540), .Z(n5543) );
  HS65_LH_CNIVX3 U8190 ( .A(n5506), .Z(n5512) );
  HS65_LH_CNIVX3 U8191 ( .A(n5541), .Z(n5525) );
  HS65_LH_AOI21X2 U8192 ( .A(n5520), .B(n5519), .C(n5518), .Z(n5523) );
  HS65_LH_CNIVX3 U8193 ( .A(n5516), .Z(n5519) );
  HS65_LH_CNIVX3 U8194 ( .A(n5517), .Z(n5518) );
  HS65_LH_CBI4I1X3 U8195 ( .A(n5531), .B(n5530), .C(n3515), .D(n5529), .Z(
        n5532) );
  HS65_LH_NAND3X2 U8196 ( .A(n5105), .B(n5104), .C(n5103), .Z(n5109) );
  HS65_LH_CBI4I1X3 U8197 ( .A(n5107), .B(n5468), .C(n5396), .D(n5106), .Z(
        n5108) );
  HS65_LH_CNIVX3 U8199 ( .A(n5302), .Z(n5296) );
  HS65_LH_CNIVX3 U8200 ( .A(n5310), .Z(n5316) );
  HS65_LH_NAND2X2 U8201 ( .A(n5327), .B(n3354), .Z(n5315) );
  HS65_LH_CNIVX3 U8202 ( .A(n5473), .Z(n5306) );
  HS65_LH_NAND2X2 U8204 ( .A(n5390), .B(n5381), .Z(n5394) );
  HS65_LH_AOI21X2 U8205 ( .A(n5386), .B(n5385), .C(n5384), .Z(n5393) );
  HS65_LH_AOI21X2 U8206 ( .A(n5391), .B(n5390), .C(n5389), .Z(n5392) );
  HS65_LH_AOI21X2 U8207 ( .A(n5403), .B(n5402), .C(n5401), .Z(n5411) );
  HS65_LH_AOI21X2 U8208 ( .A(n5409), .B(n5408), .C(n5407), .Z(n5410) );
  HS65_LH_OAI21X2 U8209 ( .A(n5397), .B(n5396), .C(n5395), .Z(n5403) );
  HS65_LH_NOR2X2 U8210 ( .A(n5379), .B(n5412), .Z(n5415) );
  HS65_LH_NAND2X2 U8211 ( .A(n5375), .B(n5402), .Z(n5379) );
  HS65_LH_NOR2X2 U8212 ( .A(n5374), .B(n5396), .Z(n5375) );
  HS65_LH_NOR2X2 U8213 ( .A(\lte_x_59/B[8] ), .B(n3360), .Z(n5374) );
  HS65_LH_AOI21X2 U8214 ( .A(n5446), .B(n5445), .C(n5444), .Z(n5455) );
  HS65_LH_AOI21X2 U8215 ( .A(n5453), .B(n5452), .C(n5451), .Z(n5454) );
  HS65_LH_OAI21X2 U8216 ( .A(n5442), .B(n3572), .C(n5502), .Z(n5445) );
  HS65_LH_NAND2X2 U8217 ( .A(n5416), .B(n5432), .Z(n5421) );
  HS65_LH_NOR2X2 U8218 ( .A(n5426), .B(n3572), .Z(n5427) );
  HS65_LH_AOI21X2 U8220 ( .A(n5347), .B(n5346), .C(n5505), .Z(n5348) );
  HS65_LH_CNIVX3 U8221 ( .A(n5471), .Z(n5358) );
  HS65_LH_AOI21X2 U8222 ( .A(n5275), .B(n5511), .C(n5355), .Z(n5359) );
  HS65_LH_NAND2X2 U8223 ( .A(n5363), .B(n5362), .Z(n5367) );
  HS65_LH_CNIVX3 U8224 ( .A(n5354), .Z(n5370) );
  HS65_LH_NOR3X1 U8225 ( .A(\sub_x_53/A[30] ), .B(n2873), .C(n5342), .Z(n4964)
         );
  HS65_LH_AOI21X2 U8226 ( .A(n4983), .B(n5582), .C(n5013), .Z(n4993) );
  HS65_LH_OAI21X2 U8227 ( .A(\sub_x_53/A[25] ), .B(n5345), .C(n4982), .Z(n4983) );
  HS65_LH_NAND3X2 U8228 ( .A(n4981), .B(n5502), .C(n5180), .Z(n4982) );
  HS65_LH_NAND3X2 U8229 ( .A(n5450), .B(n5449), .C(n5575), .Z(n4979) );
  HS65_LH_AOI21X2 U8230 ( .A(n5008), .B(n5025), .C(n5007), .Z(n5011) );
  HS65_LH_OAI21X2 U8231 ( .A(n5003), .B(n5023), .C(n5002), .Z(n5008) );
  HS65_LH_NAND2X2 U8232 ( .A(n5582), .B(n4999), .Z(n5000) );
  HS65_LH_NOR2X2 U8233 ( .A(n5500), .B(n4998), .Z(n4999) );
  HS65_LH_NOR2X2 U8234 ( .A(n3101), .B(n4997), .Z(n4998) );
  HS65_LH_OAI21X2 U8235 ( .A(n5342), .B(n5572), .C(n4229), .Z(n5014) );
  HS65_LH_NOR2X2 U8236 ( .A(n5051), .B(n5071), .Z(n5073) );
  HS65_LH_NOR2X2 U8237 ( .A(n5027), .B(n5081), .Z(n5028) );
  HS65_LH_NAND2X2 U8238 ( .A(n5026), .B(n5025), .Z(n5027) );
  HS65_LH_NOR2X2 U8239 ( .A(n5024), .B(n5023), .Z(n5026) );
  HS65_LH_AOI21X2 U8240 ( .A(n5087), .B(n5086), .C(n5085), .Z(n5112) );
  HS65_LH_NOR2X2 U8241 ( .A(n5084), .B(n5516), .Z(n5086) );
  HS65_LH_CNIVX3 U8242 ( .A(n5522), .Z(n5087) );
  HS65_LH_OAI21X2 U8243 ( .A(n5522), .B(n5517), .C(n5521), .Z(n5085) );
  HS65_LL_NOR3X1 U8244 ( .A(n5550), .B(n5384), .C(n5094), .Z(n5102) );
  HS65_LL_NAND3X2 U8245 ( .A(n5544), .B(n5545), .C(n5556), .Z(n5101) );
  HS65_LHS_XOR2X3 U8246 ( .A(\lte_x_59/B[22] ), .B(n5654), .Z(n4772) );
  HS65_LH_NOR2X2 U8247 ( .A(n5646), .B(n4526), .Z(n3784) );
  HS65_LH_NAND2X2 U8248 ( .A(n5618), .B(n5666), .Z(n3771) );
  HS65_LH_CNIVX3 U8249 ( .A(n5182), .Z(n3778) );
  HS65_LH_AOI21X2 U8250 ( .A(n9352), .B(n4997), .C(n5649), .Z(n3601) );
  HS65_LH_CNIVX3 U8251 ( .A(n4120), .Z(n3599) );
  HS65_LHS_XNOR2X3 U8252 ( .A(\sub_x_53/A[27] ), .B(n4976), .Z(n4739) );
  HS65_LHS_XNOR2X3 U8253 ( .A(n5062), .B(\lte_x_59/B[15] ), .Z(n4748) );
  HS65_LHS_XOR2X3 U8254 ( .A(n5398), .B(n2858), .Z(n4757) );
  HS65_LH_CBI4I1X3 U8255 ( .A(n3582), .B(n5231), .C(n5647), .D(n2849), .Z(
        n5236) );
  HS65_LH_AOI21X2 U8256 ( .A(n9352), .B(n5231), .C(n5649), .Z(n5237) );
  HS65_LL_NAND2AX4 U8257 ( .A(n3190), .B(n8534), .Z(n3192) );
  HS65_LHS_XNOR2X3 U8258 ( .A(n5104), .B(n5105), .Z(n4754) );
  HS65_LH_AOI21X2 U8259 ( .A(n9352), .B(n4967), .C(n5649), .Z(n3721) );
  HS65_LHS_XOR2X3 U8260 ( .A(\sub_x_53/A[23] ), .B(n4967), .Z(n4755) );
  HS65_LH_NAND2X2 U8261 ( .A(n4836), .B(n5617), .Z(n4517) );
  HS65_LL_AND2X4 U8262 ( .A(\lte_x_59/B[18] ), .B(n2864), .Z(n3908) );
  HS65_LH_NAND2X2 U8263 ( .A(n4887), .B(n4120), .Z(n4068) );
  HS65_LH_CBI4I6X2 U8264 ( .A(n9346), .B(n5376), .C(n3529), .D(n4675), .Z(
        n4067) );
  HS65_LH_AOI21X2 U8265 ( .A(n3529), .B(n3860), .C(n4682), .Z(n3861) );
  HS65_LH_NAND2X2 U8266 ( .A(n5648), .B(n5373), .Z(n3860) );
  HS65_LH_AOI21X2 U8267 ( .A(n5648), .B(n4699), .C(n5647), .Z(n4439) );
  HS65_LH_AOI21X2 U8268 ( .A(n9349), .B(n5021), .C(n4850), .Z(n4852) );
  HS65_LHS_XNOR2X3 U8269 ( .A(n5001), .B(n4984), .Z(n4742) );
  HS65_LLS_XNOR2X3 U8270 ( .A(n8764), .B(n8943), .Z(n3037) );
  HS65_LHS_XNOR2X6 U8271 ( .A(\sub_x_53/A[2] ), .B(n5088), .Z(n4769) );
  HS65_LH_AND2X4 U8272 ( .A(\u_DataPath/jaddr_i [25]), .B(
        \u_DataPath/jaddr_i [24]), .Z(n6131) );
  HS65_LH_AOI112X2 U8273 ( .A(n5648), .B(n7623), .C(n4192), .D(n3443), .Z(
        n4193) );
  HS65_LHS_XNOR2X3 U8274 ( .A(n2851), .B(n7623), .Z(n4738) );
  HS65_LH_OAI22X1 U8275 ( .A(n2854), .B(n4583), .C(n3756), .D(n4711), .Z(n3656) );
  HS65_LH_OAI22X1 U8276 ( .A(n4981), .B(n4795), .C(n5129), .D(n3101), .Z(n3657) );
  HS65_LH_CNIVX3 U8278 ( .A(n5286), .Z(n4710) );
  HS65_LH_NAND3X2 U8279 ( .A(n5270), .B(n4698), .C(n4697), .Z(n4707) );
  HS65_LH_NAND3X2 U8280 ( .A(\lte_x_59/B[18] ), .B(n5534), .C(n3371), .Z(n4698) );
  HS65_LH_OAI21X2 U8281 ( .A(n5511), .B(n4696), .C(n5432), .Z(n4697) );
  HS65_LH_NOR2X2 U8282 ( .A(n5506), .B(n3515), .Z(n4696) );
  HS65_LH_NAND3X2 U8283 ( .A(\lte_x_59/B[22] ), .B(n2869), .C(n5290), .Z(n4705) );
  HS65_LH_CBI4I1X3 U8284 ( .A(n5471), .B(n5292), .C(n5363), .D(n4703), .Z(
        n4704) );
  HS65_LH_AOI21X2 U8285 ( .A(n5286), .B(n5505), .C(n5499), .Z(n4729) );
  HS65_LH_AOI21X2 U8286 ( .A(n5503), .B(n4727), .C(n5342), .Z(n4728) );
  HS65_LH_CBI4I1X3 U8287 ( .A(n5500), .B(n5289), .C(n5012), .D(n4721), .Z(
        n4722) );
  HS65_LH_CNIVX3 U8288 ( .A(n4720), .Z(n4721) );
  HS65_LH_CNIVX3 U8289 ( .A(n5408), .Z(n4681) );
  HS65_LH_AOI21X2 U8290 ( .A(n5517), .B(n5476), .C(n5514), .Z(n4680) );
  HS65_LH_AOI21X2 U8291 ( .A(n3892), .B(n5083), .C(n4678), .Z(n4679) );
  HS65_LH_CB4I6X4 U8292 ( .A(n4687), .B(n4686), .C(n4685), .D(n4684), .Z(n4688) );
  HS65_LH_CNIVX3 U8293 ( .A(n5402), .Z(n4686) );
  HS65_LH_AOI21X2 U8294 ( .A(n5311), .B(n5335), .C(n5299), .Z(n4687) );
  HS65_LH_NAND4ABX3 U8295 ( .A(n4720), .B(n4691), .C(n5346), .D(n5572), .Z(
        n4735) );
  HS65_LH_NAND2AX4 U8296 ( .A(n4666), .B(n4659), .Z(n4670) );
  HS65_LH_NAND2X2 U8298 ( .A(n7834), .B(n5463), .Z(n5497) );
  HS65_LH_NOR3X1 U8299 ( .A(n5571), .B(n4965), .C(n4964), .Z(n4980) );
  HS65_LHS_XNOR2X3 U8300 ( .A(\sub_x_53/A[0] ), .B(n5123), .Z(n5124) );
  HS65_LH_NAND3X2 U8301 ( .A(\u_DataPath/u_idexreg/N3 ), .B(n5121), .C(n5120), 
        .Z(n5122) );
  HS65_LH_NAND2X2 U8302 ( .A(n4836), .B(n5672), .Z(n3762) );
  HS65_LH_AOI21X2 U8303 ( .A(n5648), .B(n3593), .C(n5647), .Z(n3584) );
  HS65_LH_AOI21X2 U8304 ( .A(n9352), .B(n4976), .C(n3659), .Z(n3660) );
  HS65_LH_AOI21X2 U8305 ( .A(n3529), .B(n3658), .C(n4711), .Z(n3659) );
  HS65_LH_NAND2X2 U8306 ( .A(n5648), .B(n4976), .Z(n3658) );
  HS65_LH_CNIVX3 U8307 ( .A(n4739), .Z(n3662) );
  HS65_LH_NOR2X2 U8308 ( .A(n5173), .B(n4185), .Z(n3668) );
  HS65_LH_CNIVX3 U8309 ( .A(n3751), .Z(n3631) );
  HS65_LH_CNIVX3 U8310 ( .A(n3750), .Z(n3632) );
  HS65_LH_AND2X4 U8311 ( .A(n3170), .B(n3407), .Z(n2911) );
  HS65_LH_AOI21X2 U8312 ( .A(n5965), .B(n5930), .C(n5929), .Z(n5931) );
  HS65_LH_CBI4I1X3 U8313 ( .A(n3582), .B(n5062), .C(n5647), .D(
        \lte_x_59/B[15] ), .Z(n3916) );
  HS65_LH_NAND2X2 U8314 ( .A(n4507), .B(n4942), .Z(n3915) );
  HS65_LH_AOI21X2 U8315 ( .A(n9352), .B(n5062), .C(n5649), .Z(n3917) );
  HS65_LH_OAI21X2 U8316 ( .A(n3923), .B(n5646), .C(n3922), .Z(n3924) );
  HS65_LH_NAND2X2 U8317 ( .A(n4887), .B(n4504), .Z(n3926) );
  HS65_LH_AOI21X2 U8318 ( .A(n3897), .B(n4918), .C(n3896), .Z(n3898) );
  HS65_LH_NAND2X2 U8320 ( .A(n4017), .B(n4014), .Z(n4019) );
  HS65_LH_CBI4I1X3 U8321 ( .A(n4683), .B(n5648), .C(n5647), .D(n2858), .Z(
        n4030) );
  HS65_LH_AOI21X2 U8322 ( .A(n9349), .B(n4683), .C(n4028), .Z(n4029) );
  HS65_LH_NAND2X2 U8323 ( .A(n5261), .B(n5257), .Z(n5263) );
  HS65_LH_CNIVX3 U8324 ( .A(n4494), .Z(n4495) );
  HS65_LH_CBI4I1X3 U8325 ( .A(n5648), .B(n5104), .C(n5647), .D(n3474), .Z(
        n3970) );
  HS65_LH_CNIVX3 U8326 ( .A(n5660), .Z(n3966) );
  HS65_LH_CNIVX3 U8327 ( .A(n4950), .Z(n3962) );
  HS65_LH_CNIVX3 U8328 ( .A(n4755), .Z(n3725) );
  HS65_LH_AOI21X2 U8329 ( .A(n3710), .B(n5615), .C(n3709), .Z(n3711) );
  HS65_LH_CNIVX3 U8330 ( .A(n4608), .Z(n3710) );
  HS65_LH_CNIVX3 U8331 ( .A(n5606), .Z(n3735) );
  HS65_LH_CNIVX3 U8333 ( .A(n5632), .Z(n3701) );
  HS65_LHS_XNOR2X3 U8334 ( .A(n4671), .B(n5048), .Z(n4750) );
  HS65_LH_CNIVX3 U8335 ( .A(n4625), .Z(n4626) );
  HS65_LH_CNIVX3 U8336 ( .A(n4640), .Z(n4642) );
  HS65_LH_AOI21X2 U8337 ( .A(n4581), .B(n4341), .C(n5249), .Z(n4342) );
  HS65_LL_AOI21X2 U8338 ( .A(n9349), .B(n5422), .C(n5649), .Z(n4352) );
  HS65_LHS_XOR2X3 U8340 ( .A(\sub_x_53/A[29] ), .B(n5422), .Z(n4765) );
  HS65_LH_AOI21X2 U8341 ( .A(n5618), .B(n4394), .C(n4358), .Z(n4359) );
  HS65_LH_CNIVX3 U8342 ( .A(n4356), .Z(n4357) );
  HS65_LH_NAND2X2 U8343 ( .A(n5194), .B(n4335), .Z(n4337) );
  HS65_LH_AOI21X2 U8344 ( .A(n5659), .B(n4892), .C(n4397), .Z(n4398) );
  HS65_LH_AOI21X2 U8345 ( .A(n9349), .B(n5418), .C(n5649), .Z(n4395) );
  HS65_LH_NAND2X2 U8346 ( .A(n5229), .B(n4394), .Z(n4399) );
  HS65_LH_NAND2X2 U8347 ( .A(n5661), .B(n4393), .Z(n4400) );
  HS65_LH_CNIVX3 U8348 ( .A(n4105), .Z(n4106) );
  HS65_LH_AOI21X2 U8350 ( .A(n9349), .B(n5040), .C(n4115), .Z(n4116) );
  HS65_LHS_XNOR2X3 U8352 ( .A(\lte_x_59/B[5] ), .B(n5040), .Z(n4753) );
  HS65_LH_AND2X4 U8353 ( .A(n4714), .B(n8506), .Z(n3227) );
  HS65_LH_CNIVX3 U8354 ( .A(n4902), .Z(n4903) );
  HS65_LH_CNIVX3 U8355 ( .A(n3823), .Z(n3436) );
  HS65_LH_OAI21X2 U8356 ( .A(n5004), .B(n2856), .C(n3819), .Z(n3433) );
  HS65_LH_AOI21X2 U8357 ( .A(n5648), .B(n5654), .C(n5647), .Z(n5653) );
  HS65_LH_NAND2X2 U8358 ( .A(n5608), .B(n2867), .Z(n5611) );
  HS65_LH_AOI21X2 U8359 ( .A(n5139), .B(n5618), .C(n3879), .Z(n3880) );
  HS65_LH_AOI21X2 U8360 ( .A(n9352), .B(n5373), .C(n3861), .Z(n3866) );
  HS65_LH_AOI21X2 U8362 ( .A(n5234), .B(n4441), .C(n4440), .Z(n4442) );
  HS65_LH_AOI21X2 U8363 ( .A(n5207), .B(n4892), .C(n3537), .Z(n3538) );
  HS65_LH_CNIVX3 U8365 ( .A(n4542), .Z(n4543) );
  HS65_LH_CBI4I6X2 U8366 ( .A(n9346), .B(n3415), .C(n3529), .D(n5130), .Z(
        n4549) );
  HS65_LH_CNIVX3 U8367 ( .A(n4630), .Z(n4158) );
  HS65_LHS_XNOR2X3 U8368 ( .A(\lte_x_59/B[6] ), .B(n2865), .Z(n4764) );
  HS65_LH_CNIVX3 U8369 ( .A(n3955), .Z(n3960) );
  HS65_LLS_XNOR2X3 U8370 ( .A(n2947), .B(n8762), .Z(n2959) );
  HS65_LH_CNIVX3 U8371 ( .A(n2957), .Z(n2958) );
  HS65_LH_NOR2X6 U8372 ( .A(n9236), .B(n2982), .Z(n7639) );
  HS65_LH_AOI21X2 U8374 ( .A(n9352), .B(n7623), .C(n4194), .Z(n4195) );
  HS65_LH_AOI21X2 U8375 ( .A(n4182), .B(n4181), .C(n5646), .Z(n4183) );
  HS65_LH_AOI21X2 U8376 ( .A(\lte_x_59/B[28] ), .B(n2864), .C(n4507), .Z(n4181) );
  HS65_LH_AOI21X2 U8379 ( .A(n4211), .B(n4291), .C(n4218), .Z(n4219) );
  HS65_LHS_XNOR2X3 U8380 ( .A(n8942), .B(\u_DataPath/jaddr_i [16]), .Z(n7103)
         );
  HS65_LH_AOI21X2 U8381 ( .A(n5229), .B(n4892), .C(n4801), .Z(n4802) );
  HS65_LH_AOI21X2 U8382 ( .A(n5648), .B(n4805), .C(n4804), .Z(n4812) );
  HS65_LH_OAI21X2 U8383 ( .A(n4796), .B(n4795), .C(n4794), .Z(n4797) );
  HS65_LH_CNIVX3 U8384 ( .A(n4333), .Z(n3130) );
  HS65_LL_NOR2AX3 U8385 ( .A(n2904), .B(n4735), .Z(n4692) );
  HS65_LH_NOR2X2 U8386 ( .A(n5491), .B(\u_DataPath/cw_to_ex_i [4]), .Z(n5121)
         );
  HS65_LL_AOI21X2 U8388 ( .A(n5192), .B(n5195), .C(n3576), .Z(n3577) );
  HS65_LH_NOR2X6 U8389 ( .A(n9078), .B(n9031), .Z(n7343) );
  HS65_LH_CNIVX3 U8390 ( .A(n4913), .Z(n4914) );
  HS65_LH_AOI21X2 U8392 ( .A(n4919), .B(n4918), .C(n4917), .Z(n4920) );
  HS65_LL_NOR3AX2 U8393 ( .A(n3926), .B(n3925), .C(n3924), .Z(n3927) );
  HS65_LH_AOI21X2 U8394 ( .A(n5234), .B(n3919), .C(n3918), .Z(n3928) );
  HS65_LH_AOI21X2 U8395 ( .A(n4951), .B(n4616), .C(n3906), .Z(n3931) );
  HS65_LH_CNIVX3 U8396 ( .A(n4011), .Z(n4012) );
  HS65_LH_CNIVX3 U8397 ( .A(n4570), .Z(n4571) );
  HS65_LH_AOI21X2 U8398 ( .A(n4508), .B(n4507), .C(n4506), .Z(n4509) );
  HS65_LH_CNIVX3 U8400 ( .A(n4938), .Z(n4492) );
  HS65_LH_AND2X4 U8401 ( .A(n5405), .B(n4051), .Z(n2906) );
  HS65_LH_CNIVX3 U8404 ( .A(n4771), .Z(n4613) );
  HS65_LH_AOI21X2 U8405 ( .A(n9352), .B(n5030), .C(n4610), .Z(n4611) );
  HS65_LH_OAI22X1 U8406 ( .A(n4954), .B(n3913), .C(n4609), .D(n5646), .Z(n4621) );
  HS65_LH_OAI21X2 U8407 ( .A(n4113), .B(n5201), .C(n4065), .Z(n4075) );
  HS65_LH_AOI21X2 U8409 ( .A(n5618), .B(n5203), .C(n5202), .Z(n5220) );
  HS65_LH_OAI21X2 U8410 ( .A(n3382), .B(n5179), .C(n5178), .Z(n5185) );
  HS65_LH_NAND2X2 U8412 ( .A(n4516), .B(n4491), .Z(n4161) );
  HS65_LHS_XOR2X3 U8413 ( .A(n3856), .B(n4929), .Z(n3888) );
  HS65_LH_CNIVX3 U8414 ( .A(n4880), .Z(n3855) );
  HS65_LH_NAND2X2 U8415 ( .A(n4836), .B(n4835), .Z(n4837) );
  HS65_LH_CNIVX3 U8416 ( .A(n4575), .Z(n4539) );
  HS65_LH_AOI21X2 U8417 ( .A(n4546), .B(n4545), .C(n5201), .Z(n4547) );
  HS65_LH_CNIVX3 U8418 ( .A(n4541), .Z(n4546) );
  HS65_LH_AOI21X2 U8419 ( .A(\lte_x_59/B[4] ), .B(n4544), .C(n4543), .Z(n4545)
         );
  HS65_LH_NOR2AX3 U8420 ( .A(n4557), .B(n4556), .Z(n4566) );
  HS65_LH_AOI21X2 U8421 ( .A(n9352), .B(n5088), .C(n4549), .Z(n4557) );
  HS65_LH_CNIVX3 U8422 ( .A(n4643), .Z(n4142) );
  HS65_LH_IVX9 U8423 ( .A(n3409), .Z(n3237) );
  HS65_LH_NOR2X2 U8424 ( .A(n9084), .B(n9082), .Z(n7693) );
  HS65_LH_AOI21X2 U8425 ( .A(n9082), .B(n7734), .C(n7690), .Z(n7692) );
  HS65_LH_NAND2X2 U8427 ( .A(n4836), .B(n5243), .Z(n4177) );
  HS65_LH_AOI21X2 U8428 ( .A(n5661), .B(n5228), .C(n4186), .Z(n4201) );
  HS65_LH_AOI21X2 U8430 ( .A(n5234), .B(n4199), .C(n4198), .Z(n4200) );
  HS65_LH_NAND2X2 U8431 ( .A(n2851), .B(n7623), .Z(n4206) );
  HS65_LH_IVX9 U8432 ( .A(n8683), .Z(n7742) );
  HS65_LH_IVX9 U8433 ( .A(n8695), .Z(n7753) );
  HS65_LH_IVX9 U8434 ( .A(n8694), .Z(n3123) );
  HS65_LH_IVX9 U8435 ( .A(n8699), .Z(n3125) );
  HS65_LH_IVX9 U8437 ( .A(n8709), .Z(n3124) );
  HS65_LH_IVX9 U8438 ( .A(n8705), .Z(n7769) );
  HS65_LH_IVX9 U8439 ( .A(n8708), .Z(n7756) );
  HS65_LH_IVX9 U8440 ( .A(n8706), .Z(n7766) );
  HS65_LH_IVX9 U8441 ( .A(n8711), .Z(n3121) );
  HS65_LH_IVX9 U8442 ( .A(n8701), .Z(n3119) );
  HS65_LH_IVX9 U8443 ( .A(n8707), .Z(n3118) );
  HS65_LH_IVX9 U8444 ( .A(n8710), .Z(n7705) );
  HS65_LH_IVX9 U8445 ( .A(n8712), .Z(n7785) );
  HS65_LH_NOR3X1 U8446 ( .A(n7636), .B(n7778), .C(n7772), .Z(n7309) );
  HS65_LH_CBI4I1X3 U8447 ( .A(n8116), .B(n7698), .C(n7689), .D(n7697), .Z(
        n8118) );
  HS65_LH_OAI22X1 U8448 ( .A(n7738), .B(n7690), .C(n9084), .D(n7688), .Z(n7689) );
  HS65_LL_AND2X4 U8449 ( .A(n5682), .B(n5681), .Z(n5685) );
  HS65_LL_NOR3AX2 U8450 ( .A(n7873), .B(n5680), .C(n5679), .Z(n5682) );
  HS65_LLS_XNOR2X3 U8451 ( .A(n3393), .B(n3392), .Z(n3514) );
  HS65_LLS_XNOR2X3 U8452 ( .A(n3638), .B(n3637), .Z(n3697) );
  HS65_LH_IVX2 U8453 ( .A(n7622), .Z(n7621) );
  HS65_LH_NAND3X2 U8454 ( .A(n7089), .B(n9031), .C(n9078), .Z(n8145) );
  HS65_LH_NAND3X5 U8455 ( .A(n3011), .B(n9078), .C(n2946), .Z(n8147) );
  HS65_LH_IVX9 U8456 ( .A(n7840), .Z(n8608) );
  HS65_LH_OAI21X2 U8457 ( .A(n9084), .B(n7775), .C(n7774), .Z(n7779) );
  HS65_LH_CNIVX3 U8459 ( .A(n6066), .Z(n6009) );
  HS65_LH_CNIVX3 U8461 ( .A(n5947), .Z(n5948) );
  HS65_LH_CNIVX3 U8463 ( .A(n8258), .Z(n3241) );
  HS65_LH_CNIVX3 U8464 ( .A(n6061), .Z(n6062) );
  HS65_LH_CNIVX3 U8465 ( .A(n5952), .Z(n5953) );
  HS65_LH_AOI22X1 U8466 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][27] ), .Z(n7460)
         );
  HS65_LH_AO22X4 U8467 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][27] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ), .Z(n7463)
         );
  HS65_LH_AO22X4 U8468 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][27] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ), .Z(n7462)
         );
  HS65_LH_AOI22X1 U8469 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][27] ), .Z(n7461)
         );
  HS65_LH_AOI22X1 U8470 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][27] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][27] ), .D(n6746), 
        .Z(n7459) );
  HS65_LH_AO22X4 U8471 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][27] ), .D(
        n6675), .Z(n7457) );
  HS65_LH_AO22X4 U8472 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][27] ), .B(n7578), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ), .Z(n7453)
         );
  HS65_LH_AOI22X1 U8473 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][27] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][27] ), .D(n2890), 
        .Z(n7454) );
  HS65_LH_AO22X4 U8475 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ), .D(
        n6627), .Z(n6310) );
  HS65_LH_AO22X4 U8476 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][14] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ), .D(
        n6629), .Z(n6309) );
  HS65_LH_AO22X4 U8477 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][14] ), .D(
        n7292), .Z(n6320) );
  HS65_LH_AOI22X1 U8478 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ), .D(
        n7296), .Z(n6318) );
  HS65_LH_AO22X4 U8479 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][14] ), .D(
        n6382), .Z(n6321) );
  HS65_LH_AO22X4 U8480 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][14] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][14] ), .D(
        n6635), .Z(n6316) );
  HS65_LH_AO22X4 U8481 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][14] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][14] ), .D(
        n6619), .Z(n6305) );
  HS65_LH_AO22X4 U8482 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][14] ), .D(
        n9371), .Z(n6306) );
  HS65_LH_AOI22X1 U8483 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][14] ), .D(
        n6363), .Z(n6307) );
  HS65_LH_AO22X4 U8484 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][14] ), .D(
        n7586), .Z(n7371) );
  HS65_LH_AO22X4 U8485 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][14] ), .D(
        n6675), .Z(n7372) );
  HS65_LH_AOI22X1 U8486 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][14] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ), .Z(n7380)
         );
  HS65_LH_AOI22X1 U8487 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][14] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ), .Z(n7379)
         );
  HS65_LH_AOI22X1 U8488 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][14] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][14] ), .D(n6740), 
        .Z(n7369) );
  HS65_LH_AOI22X1 U8489 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][14] ), .Z(n7375)
         );
  HS65_LH_AO22X4 U8490 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ), .D(
        n7319), .Z(n7188) );
  HS65_LH_AOI22X1 U8491 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ), .D(
        n6670), .Z(n7187) );
  HS65_LH_AOI22X1 U8492 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][15] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ), .D(n6740), 
        .Z(n7186) );
  HS65_LH_AO22X4 U8493 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ), .B(n9373), 
        .C(n7311), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ), .Z(n7184)
         );
  HS65_LH_AO22X4 U8494 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][15] ), .Z(n7198)
         );
  HS65_LH_AO22X4 U8495 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][15] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][15] ), .Z(n7199)
         );
  HS65_LH_AOI22X1 U8496 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][15] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][15] ), .Z(n7192)
         );
  HS65_LH_AO22X4 U8497 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][11] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][11] ), .Z(n7067)
         );
  HS65_LH_AOI22X1 U8498 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][11] ), .Z(n7065)
         );
  HS65_LH_AOI22X1 U8499 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][11] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ), .D(
        n6670), .Z(n7059) );
  HS65_LH_AOI22X1 U8500 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][11] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][11] ), .D(n2890), 
        .Z(n7058) );
  HS65_LH_AOI22X1 U8501 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][11] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][11] ), .D(n6746), 
        .Z(n7063) );
  HS65_LH_CNIVX3 U8502 ( .A(n9232), .Z(n4005) );
  HS65_LH_AOI22X1 U8503 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][19] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ), .D(n6746), 
        .Z(n6751) );
  HS65_LH_AOI22X1 U8504 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][19] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ), .D(
        n6670), .Z(n6744) );
  HS65_LH_AOI22X1 U8505 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][19] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][19] ), .D(n2890), 
        .Z(n6743) );
  HS65_LH_AO22X4 U8506 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][19] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][19] ), .Z(n6758)
         );
  HS65_LH_CNIVX3 U8507 ( .A(n9218), .Z(n5702) );
  HS65_LH_AO22X4 U8509 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ), .D(
        n7586), .Z(n7391) );
  HS65_LH_AO22X4 U8510 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][3] ), .D(n6675), .Z(n7392) );
  HS65_LH_AOI22X1 U8511 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][3] ), .Z(n7400)
         );
  HS65_LH_AOI22X1 U8512 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][3] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][3] ), .Z(n7399)
         );
  HS65_LH_AOI22X1 U8513 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][3] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][3] ), .Z(n7396)
         );
  HS65_LH_AOI22X1 U8514 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][10] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][10] ), .D(n6740), 
        .Z(n7206) );
  HS65_LH_AO22X4 U8515 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][10] ), .B(n7578), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ), .Z(n7205)
         );
  HS65_LH_AO22X4 U8516 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ), .B(n9373), 
        .C(n7311), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ), .Z(n7204)
         );
  HS65_LH_AOI22X1 U8517 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][10] ), .Z(n7217)
         );
  HS65_LH_AOI22X1 U8518 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][10] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][10] ), .Z(n7216)
         );
  HS65_LH_AO22X4 U8519 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][10] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][10] ), .Z(n7219)
         );
  HS65_LH_AO22X4 U8520 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][10] ), .Z(n7218)
         );
  HS65_LH_AOI22X1 U8521 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][10] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][10] ), .Z(n7212)
         );
  HS65_LH_AO22X4 U8522 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][10] ), .D(
        n7319), .Z(n7208) );
  HS65_LH_AOI22X1 U8523 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][23] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][23] ), .D(n6740), 
        .Z(n7226) );
  HS65_LH_AO22X4 U8524 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][23] ), .B(n7429), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ), .Z(n7225)
         );
  HS65_LH_AO22X4 U8525 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][23] ), .B(n9373), 
        .C(n7311), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][23] ), .Z(n7224)
         );
  HS65_LH_AOI22X1 U8526 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ), .Z(n7237)
         );
  HS65_LH_AOI22X1 U8527 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][23] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][23] ), .Z(n7236)
         );
  HS65_LH_AO22X4 U8528 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][23] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][23] ), .Z(n7239)
         );
  HS65_LH_AO22X4 U8529 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][23] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][23] ), .Z(n7238)
         );
  HS65_LH_AOI22X1 U8530 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][23] ), .Z(n7232)
         );
  HS65_LH_AO22X4 U8531 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][23] ), .D(
        n7319), .Z(n7228) );
  HS65_LH_AO22X4 U8532 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][30] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ), .D(
        n6627), .Z(n6135) );
  HS65_LH_AO22X4 U8533 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][30] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ), .D(
        n6629), .Z(n6134) );
  HS65_LH_AO22X4 U8534 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ), .D(
        n7292), .Z(n6156) );
  HS65_LH_AOI22X1 U8535 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][30] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ), .D(
        n7296), .Z(n6154) );
  HS65_LH_AO22X4 U8536 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][30] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ), .D(
        n6382), .Z(n6157) );
  HS65_LH_AO22X4 U8537 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ), .D(
        n6637), .Z(n6143) );
  HS65_LH_AO22X4 U8538 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ), .D(
        n6635), .Z(n6144) );
  HS65_LH_AO22X4 U8539 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ), .D(
        n6619), .Z(n6127) );
  HS65_LH_AO22X4 U8540 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][30] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ), .D(
        n9371), .Z(n6128) );
  HS65_LH_AOI22X1 U8541 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][30] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][30] ), .D(n6746), 
        .Z(n7413) );
  HS65_LH_AO22X4 U8542 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][30] ), .B(n6747), 
        .C(n6675), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][30] ), .Z(n7412)
         );
  HS65_LH_AO22X4 U8543 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][30] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ), .Z(n7408)
         );
  HS65_LH_AO22X4 U8544 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][30] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][30] ), .Z(n7407)
         );
  HS65_LH_AOI22X1 U8545 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][30] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][30] ), .Z(n7421)
         );
  HS65_LH_AO22X4 U8546 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][30] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][30] ), .Z(n7423)
         );
  HS65_LH_AO22X4 U8547 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ), .B(n7578), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][30] ), .D(
        n6952), .Z(n7419) );
  HS65_LH_AOI22X1 U8548 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][30] ), .D(n2890), 
        .Z(n7416) );
  HS65_LH_AND2X4 U8549 ( .A(n5450), .B(n4303), .Z(n2915) );
  HS65_LH_AO22X4 U8550 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][12] ), .D(
        n7319), .Z(n6791) );
  HS65_LH_AOI22X1 U8551 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][12] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ), .D(
        n6670), .Z(n6790) );
  HS65_LH_AOI22X1 U8552 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][12] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][12] ), .D(n6740), 
        .Z(n6789) );
  HS65_LH_AO22X4 U8553 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][12] ), .B(n7429), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ), .Z(n6788)
         );
  HS65_LH_AO22X4 U8554 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ), .B(n9373), 
        .C(n7311), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ), .Z(n6787)
         );
  HS65_LH_AO22X4 U8555 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][12] ), .Z(n6801)
         );
  HS65_LH_AO22X4 U8556 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][12] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][12] ), .Z(n6802)
         );
  HS65_LH_AOI22X1 U8557 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][12] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][12] ), .Z(n6795)
         );
  HS65_LH_AO22X4 U8558 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][7] ), .D(
        n7319), .Z(n6723) );
  HS65_LH_AOI22X1 U8559 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][7] ), .Z(n6732)
         );
  HS65_LH_AOI22X1 U8560 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][7] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][7] ), .Z(n6731)
         );
  HS65_LH_AO22X4 U8561 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][7] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ), .Z(n6734)
         );
  HS65_LH_AO22X4 U8562 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][7] ), .Z(n6733)
         );
  HS65_LH_AOI22X1 U8563 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][7] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][7] ), .Z(n6727)
         );
  HS65_LH_AO22X4 U8564 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ), .B(n9373), 
        .C(n7311), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ), .Z(n6719) );
  HS65_LH_AO22X4 U8565 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][7] ), .B(n7429), 
        .C(n6952), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ), .Z(n6720) );
  HS65_LH_AOI22X1 U8566 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][7] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][7] ), .D(n6740), 
        .Z(n6721) );
  HS65_LH_AOI22X1 U8567 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][13] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ), .D(
        n6625), .Z(n7168) );
  HS65_LH_AO22X4 U8568 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][13] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ), .D(
        n6627), .Z(n7167) );
  HS65_LH_AO22X4 U8569 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][13] ), .D(
        n6382), .Z(n7179) );
  HS65_LH_AOI22X1 U8570 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ), .D(
        n7296), .Z(n7176) );
  HS65_LH_AO22X4 U8571 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ), .D(
        n6635), .Z(n7175) );
  HS65_LH_AO22X4 U8572 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][13] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ), .D(
        n6619), .Z(n7161) );
  HS65_LH_AO22X4 U8573 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ), .D(
        n9372), .Z(n7162) );
  HS65_LH_AO22X4 U8574 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][13] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ), .Z(n6987)
         );
  HS65_LH_AOI22X1 U8575 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][13] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][13] ), .Z(n6985)
         );
  HS65_LH_AOI22X1 U8576 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][13] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][13] ), .D(
        n6670), .Z(n6979) );
  HS65_LH_AOI22X1 U8577 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][13] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][13] ), .D(n2890), 
        .Z(n6978) );
  HS65_LH_AOI22X1 U8578 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][13] ), .D(n6746), 
        .Z(n6983) );
  HS65_LH_AOI22X1 U8579 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][29] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ), .Z(n7527)
         );
  HS65_LH_AOI22X1 U8580 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][29] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][29] ), .Z(n7526)
         );
  HS65_LH_AO22X4 U8581 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][29] ), .D(
        n7586), .Z(n7518) );
  HS65_LH_AO22X4 U8582 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][29] ), .D(
        n6675), .Z(n7519) );
  HS65_LH_AOI22X1 U8583 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][29] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][29] ), .D(n6740), 
        .Z(n7514) );
  HS65_LH_AO22X4 U8584 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][21] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][21] ), .D(
        n6627), .Z(n6190) );
  HS65_LH_AO22X4 U8585 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][21] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][21] ), .D(
        n6629), .Z(n6189) );
  HS65_LH_AO22X4 U8586 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ), .D(
        n7292), .Z(n6199) );
  HS65_LH_AOI22X1 U8587 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ), .D(
        n7296), .Z(n6197) );
  HS65_LH_AO22X4 U8588 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][21] ), .D(
        n6382), .Z(n6200) );
  HS65_LH_AOI22X1 U8589 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][21] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ), .D(
        n6171), .Z(n6194) );
  HS65_LH_AO22X4 U8590 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ), .D(
        n6635), .Z(n6196) );
  HS65_LH_AO22X4 U8591 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][21] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ), .D(
        n6619), .Z(n6185) );
  HS65_LH_AO22X4 U8592 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ), .D(
        n9372), .Z(n6186) );
  HS65_LH_AOI22X1 U8593 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ), .D(
        n6363), .Z(n6187) );
  HS65_LH_AOI22X1 U8594 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][21] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][21] ), .D(
        n2891), .Z(n7584) );
  HS65_LH_AOI22X1 U8595 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][21] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][21] ), .D(n2890), 
        .Z(n7583) );
  HS65_LH_AO22X4 U8596 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][21] ), .B(n7578), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][21] ), .Z(n7582)
         );
  HS65_LH_AOI22X1 U8597 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][21] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][21] ), .D(n6746), 
        .Z(n7591) );
  HS65_LH_AO22X4 U8598 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][21] ), .D(
        n6675), .Z(n7589) );
  HS65_LH_AOI22X1 U8599 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][21] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][21] ), .Z(n7596)
         );
  HS65_LH_AO22X4 U8600 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ), .Z(n7597)
         );
  HS65_LH_AO22X4 U8601 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][21] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ), .Z(n7598)
         );
  HS65_LH_AOI22X1 U8602 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][5] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][5] ), .D(n6740), 
        .Z(n6701) );
  HS65_LH_AO22X4 U8603 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][5] ), .B(n7429), 
        .C(n6952), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ), .Z(n6700) );
  HS65_LH_AO22X4 U8604 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ), .B(n9373), 
        .C(n7311), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][5] ), .Z(n6699) );
  HS65_LH_AOI22X1 U8605 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][5] ), .Z(n6712)
         );
  HS65_LH_AOI22X1 U8606 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][5] ), .Z(n6711)
         );
  HS65_LH_AO22X4 U8607 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][5] ), .Z(n6714)
         );
  HS65_LH_AO22X4 U8608 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][5] ), .Z(n6713)
         );
  HS65_LH_AOI22X1 U8609 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][5] ), .Z(n6707)
         );
  HS65_LH_AO22X4 U8610 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][5] ), .D(
        n7319), .Z(n6703) );
  HS65_LH_AO22X4 U8611 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][25] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][25] ), .Z(n7047)
         );
  HS65_LH_AOI22X1 U8612 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][25] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][25] ), .Z(n7045)
         );
  HS65_LH_AOI22X1 U8613 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][25] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ), .D(
        n6670), .Z(n7039) );
  HS65_LH_AOI22X1 U8614 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][25] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][25] ), .D(n2890), 
        .Z(n7038) );
  HS65_LH_AOI22X1 U8615 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][25] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][25] ), .D(n6746), 
        .Z(n7043) );
  HS65_LH_AO22X4 U8616 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][9] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][9] ), .Z(n7027)
         );
  HS65_LH_AOI22X1 U8617 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][9] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][9] ), .Z(n7025)
         );
  HS65_LH_AOI22X1 U8618 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][9] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ), .D(
        n6670), .Z(n7019) );
  HS65_LH_AOI22X1 U8619 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][9] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][9] ), .D(n2890), 
        .Z(n7018) );
  HS65_LH_AOI22X1 U8620 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][9] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][9] ), .D(n6746), 
        .Z(n7023) );
  HS65_LH_AO22X4 U8621 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][24] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][24] ), .D(
        n6627), .Z(n6290) );
  HS65_LH_AO22X4 U8622 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][24] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][24] ), .D(
        n6629), .Z(n6289) );
  HS65_LH_AOI22X1 U8623 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][24] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ), .D(
        n7296), .Z(n6297) );
  HS65_LH_AO22X4 U8624 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][24] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][24] ), .D(
        n6382), .Z(n6300) );
  HS65_LH_AO22X4 U8625 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ), .D(
        n6637), .Z(n6295) );
  HS65_LH_AO22X4 U8626 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ), .D(
        n6635), .Z(n6296) );
  HS65_LH_AO22X4 U8627 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][24] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ), .D(
        n6619), .Z(n6285) );
  HS65_LH_AO22X4 U8628 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][24] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ), .D(
        n9371), .Z(n6286) );
  HS65_LH_AO22X4 U8629 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][24] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][24] ), .Z(n7569)
         );
  HS65_LH_AO22X4 U8630 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][24] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ), .Z(n7568)
         );
  HS65_LH_AOI22X1 U8631 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][24] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][24] ), .Z(n7567)
         );
  HS65_LH_AOI22X1 U8632 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][24] ), .D(n6746), 
        .Z(n7565) );
  HS65_LH_AO22X4 U8633 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ), .D(
        n6675), .Z(n7563) );
  HS65_LH_AO22X4 U8634 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][24] ), .B(n7578), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][24] ), .Z(n7559)
         );
  HS65_LH_AOI22X1 U8635 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][24] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][24] ), .D(n2890), 
        .Z(n7560) );
  HS65_LH_AO22X4 U8636 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][28] ), .D(
        n7586), .Z(n7496) );
  HS65_LH_AO22X4 U8637 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ), .D(
        n6675), .Z(n7497) );
  HS65_LH_AOI22X1 U8638 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][28] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][28] ), .Z(n7501)
         );
  HS65_LH_AO22X4 U8639 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][22] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][22] ), .D(
        n6627), .Z(n6270) );
  HS65_LH_AO22X4 U8640 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][22] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][22] ), .D(
        n6629), .Z(n6269) );
  HS65_LH_AOI22X1 U8641 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ), .B(n6385), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ), .D(
        n7296), .Z(n6277) );
  HS65_LH_AO22X4 U8642 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ), .D(
        n6382), .Z(n6280) );
  HS65_LH_AO22X4 U8643 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ), .D(
        n6637), .Z(n6275) );
  HS65_LH_AO22X4 U8644 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ), .B(n6634), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ), .D(
        n6635), .Z(n6276) );
  HS65_LH_AO22X4 U8645 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ), .D(
        n6619), .Z(n6265) );
  HS65_LH_AO22X4 U8646 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][22] ), .D(
        n9372), .Z(n6266) );
  HS65_LH_AO22X4 U8647 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][22] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][22] ), .Z(n7007)
         );
  HS65_LH_AOI22X1 U8648 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][22] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][22] ), .Z(n7005)
         );
  HS65_LH_AOI22X1 U8649 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][22] ), .D(
        n6670), .Z(n6999) );
  HS65_LH_AOI22X1 U8650 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][22] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][22] ), .D(n2890), 
        .Z(n6998) );
  HS65_LH_AOI22X1 U8651 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][22] ), .D(n6746), 
        .Z(n7003) );
  HS65_LH_CNIVX3 U8652 ( .A(n9213), .Z(n5697) );
  HS65_LH_AOI22X1 U8653 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ), .B(n6690), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][4] ), .Z(n7359)
         );
  HS65_LH_AOI22X1 U8654 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ), .B(n6689), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][4] ), .Z(n7360)
         );
  HS65_LH_AO22X4 U8655 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][4] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][4] ), .Z(n7358)
         );
  HS65_LH_AOI22X1 U8656 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][4] ), .B(n6753), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][4] ), .Z(n7356)
         );
  HS65_LH_AO22X4 U8657 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][4] ), .B(n6681), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][4] ), .Z(n7357)
         );
  HS65_LH_AO22X4 U8658 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][4] ), .B(n7578), 
        .C(n6952), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ), .Z(n7348) );
  HS65_LH_AOI22X1 U8659 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][4] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][4] ), .D(n2890), 
        .Z(n7349) );
  HS65_LH_AOI22X1 U8660 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][4] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ), .D(n6746), 
        .Z(n7354) );
  HS65_LH_AO22X4 U8661 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][4] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][4] ), .D(n6675), .Z(n7352) );
  HS65_LH_AO22X4 U8662 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][8] ), .D(
        n7319), .Z(n6771) );
  HS65_LH_AOI22X1 U8663 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][8] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ), .D(
        n6670), .Z(n6770) );
  HS65_LH_AOI22X1 U8664 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][8] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][8] ), .D(n6740), 
        .Z(n6769) );
  HS65_LH_AO22X4 U8665 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][8] ), .B(n7429), 
        .C(n7310), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ), .Z(n6768) );
  HS65_LH_AO22X4 U8666 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ), .B(n9373), 
        .C(n7311), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ), .Z(n6767) );
  HS65_LH_AO22X4 U8667 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ), .Z(n6781)
         );
  HS65_LH_AO22X4 U8668 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][8] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][8] ), .Z(n6782)
         );
  HS65_LH_AOI22X1 U8669 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][8] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][8] ), .Z(n6775)
         );
  HS65_LH_AOI22X1 U8670 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][20] ), .B(n7524), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][20] ), .Z(n7481)
         );
  HS65_LH_AOI22X1 U8671 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][20] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][20] ), .Z(n7480)
         );
  HS65_LH_AO22X4 U8672 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][20] ), .D(
        n7586), .Z(n7476) );
  HS65_LH_AO22X4 U8673 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][20] ), .D(
        n6675), .Z(n7477) );
  HS65_LH_AO22X4 U8674 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][20] ), .B(n7578), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ), .Z(n7473)
         );
  HS65_LH_AOI22X1 U8675 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ), .D(
        n2891), .Z(n7541) );
  HS65_LH_AOI22X1 U8676 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][16] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][16] ), .D(n2890), 
        .Z(n7540) );
  HS65_LH_AO22X4 U8677 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][16] ), .B(n7578), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ), .Z(n7539)
         );
  HS65_LH_AOI22X1 U8678 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][16] ), .D(n6746), 
        .Z(n7545) );
  HS65_LH_AO22X4 U8679 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ), .B(n6747), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ), .D(
        n6675), .Z(n7543) );
  HS65_LH_AOI22X1 U8680 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][16] ), .B(n6753), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][16] ), .Z(n7547)
         );
  HS65_LH_AO22X4 U8681 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][16] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ), .Z(n7548)
         );
  HS65_LH_AO22X4 U8682 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][16] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ), .Z(n7549)
         );
  HS65_LH_AOI22X1 U8683 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][2] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][2] ), .D(n2890), 
        .Z(n6955) );
  HS65_LH_AO22X4 U8684 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][2] ), .B(n7578), 
        .C(n6952), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ), .Z(n6954) );
  HS65_LH_AOI22X1 U8685 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ), .B(n6690), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][2] ), .Z(n6968)
         );
  HS65_LH_AOI22X1 U8686 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ), .B(n6689), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ), .Z(n6969)
         );
  HS65_LH_AOI22X1 U8687 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][2] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ), .D(n6746), 
        .Z(n6961) );
  HS65_LH_AO22X4 U8688 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][2] ), .D(
        n7586), .Z(n6958) );
  HS65_LH_AO22X4 U8689 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][2] ), .B(n6681), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][2] ), .Z(n6964)
         );
  HS65_LH_AOI22X1 U8690 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ), .B(n6753), 
        .C(n6683), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][2] ), .Z(n6963)
         );
  HS65_LH_AO22X4 U8691 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][2] ), .B(n6680), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][2] ), .Z(n6965)
         );
  HS65_LH_CNIVX3 U8692 ( .A(n4261), .Z(n4266) );
  HS65_LH_AOI22X1 U8693 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][18] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ), .D(
        n6670), .Z(n6330) );
  HS65_LH_CNIVX3 U8694 ( .A(n9220), .Z(n5700) );
  HS65_LH_AOI22X1 U8695 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ), .B(n6162), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ), .D(
        n2888), .Z(n6477) );
  HS65_LH_AOI22X1 U8696 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ), .B(n6371), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][6] ), .D(
        n7272), .Z(n6481) );
  HS65_LH_AO22X4 U8697 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ), .B(n6628), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][6] ), .D(
        n7276), .Z(n6479) );
  HS65_LH_AO22X4 U8698 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][6] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][6] ), .D(
        n6383), .Z(n6489) );
  HS65_LH_AOI22X1 U8699 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][6] ), .D(
        n6171), .Z(n6484) );
  HS65_LH_AO22X4 U8700 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ), .B(n6636), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ), .D(
        n7284), .Z(n6485) );
  HS65_LH_AO22X4 U8701 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][6] ), .D(
        n7319), .Z(n7248) );
  HS65_LH_AOI22X1 U8702 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][6] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][6] ), .D(
        n6670), .Z(n7247) );
  HS65_LH_AOI22X1 U8703 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][6] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][6] ), .D(n6740), 
        .Z(n7246) );
  HS65_LH_AO22X4 U8704 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][6] ), .B(n9373), 
        .C(n7311), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][6] ), .Z(n7244) );
  HS65_LH_AO22X4 U8705 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ), .Z(n7258)
         );
  HS65_LH_AO22X4 U8706 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][6] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][6] ), .Z(n7259)
         );
  HS65_LH_AOI22X1 U8707 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][6] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][6] ), .Z(n7252)
         );
  HS65_LH_AO22X4 U8708 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][0] ), .D(
        n7586), .Z(n7435) );
  HS65_LH_AO22X4 U8709 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][0] ), .D(n6675), .Z(n7436) );
  HS65_LH_AOI22X1 U8710 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][0] ), .B(n6951), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ), .D(
        n6670), .Z(n7433) );
  HS65_LH_AOI22X1 U8711 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][0] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ), .Z(n7440)
         );
  HS65_LH_CNIVX3 U8712 ( .A(n7638), .Z(n7641) );
  HS65_LH_NAND2X2 U8713 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .B(
        \u_DataPath/immediate_ext_dec_i [0]), .Z(n8089) );
  HS65_LH_AO22X4 U8714 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ), .B(n7320), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ), .D(
        n7319), .Z(n6676) );
  HS65_LH_AOI22X1 U8715 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ), .B(n6689), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ), .Z(n6692)
         );
  HS65_LH_AOI22X1 U8716 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ), .B(n6690), 
        .C(n6967), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ), .Z(n6691)
         );
  HS65_LH_AO22X4 U8717 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ), .B(n7330), 
        .C(n7329), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ), .Z(n6694)
         );
  HS65_LH_AO22X4 U8718 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ), .B(n7332), 
        .C(n7331), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ), .Z(n6693)
         );
  HS65_LH_AOI22X1 U8719 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][31] ), .B(n7525), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][31] ), .Z(n6685)
         );
  HS65_LH_AO22X4 U8720 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ), .B(n9373), 
        .C(n7311), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][31] ), .Z(n6671)
         );
  HS65_LH_AO22X4 U8721 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][31] ), .B(n7429), 
        .C(n6952), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ), .Z(n6672)
         );
  HS65_LH_AOI22X1 U8722 ( .A(n7428), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][31] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][31] ), .D(n6740), 
        .Z(n6673) );
  HS65_LHS_XOR2X3 U8723 ( .A(n7742), .B(n7741), .Z(\u_DataPath/pc_4_i [6]) );
  HS65_LHS_XOR2X3 U8724 ( .A(n7758), .B(n7757), .Z(\u_DataPath/pc_4_i [18]) );
  HS65_LH_BFX9 U8725 ( .A(n8288), .Z(n7897) );
  HS65_LH_CNIVX3 U8726 ( .A(n8117), .Z(n8058) );
  HS65_LH_OR2X4 U8727 ( .A(n8911), .B(n9202), .Z(n5919) );
  HS65_LH_IVX2 U8728 ( .A(Data_out_fromRAM[31]), .Z(n8420) );
  HS65_LH_IVX44 U8736 ( .A(n8270), .Z(nibble[0]) );
  HS65_LH_IVX40 U8737 ( .A(\u_DataPath/pc_4_i [2]), .Z(addr_to_iram[0]) );
  HS65_LH_IVX40 U8738 ( .A(n7669), .Z(addr_to_iram[2]) );
  HS65_LH_IVX40 U8739 ( .A(n7745), .Z(addr_to_iram[3]) );
  HS65_LH_IVX40 U8740 ( .A(n7667), .Z(addr_to_iram[5]) );
  HS65_LH_IVX40 U8741 ( .A(n7769), .Z(addr_to_iram[19]) );
  HS65_LH_IVX40 U8742 ( .A(n7756), .Z(addr_to_iram[20]) );
  HS65_LH_IVX40 U8743 ( .A(n7766), .Z(addr_to_iram[21]) );
  HS65_LH_IVX40 U8744 ( .A(n7705), .Z(addr_to_iram[27]) );
  HS65_LH_NAND2AX4 U8745 ( .A(n8480), .B(n9110), .Z(n8048) );
  HS65_LH_AO22X4 U8746 ( .A(n9185), .B(n8067), .C(n8966), .D(n8066), .Z(
        \u_DataPath/RFaddr_out_memwb_i [1]) );
  HS65_LH_AO22X4 U8747 ( .A(n8765), .B(n9252), .C(n9325), .D(n9153), .Z(
        \u_DataPath/jaddr_i [22]) );
  HS65_LH_NAND2AX4 U8748 ( .A(n8480), .B(\u_DataPath/cw_exmem_i [10]), .Z(
        n7833) );
  HS65_LH_CNIVX3 U8749 ( .A(n8761), .Z(n8063) );
  HS65_LH_CNIVX3 U8750 ( .A(n8764), .Z(n8065) );
  HS65_LH_NOR2X2 U8751 ( .A(n8177), .B(rst), .Z(n8580) );
  HS65_LH_NAND2AX4 U8752 ( .A(n8480), .B(n9238), .Z(n8137) );
  HS65_LH_AO222X4 U8753 ( .A(n7896), .B(\u_DataPath/pc_4_i [26]), .C(n7893), 
        .D(\u_DataPath/jump_address_i [26]), .E(n8940), .F(n7887), .Z(n8646)
         );
  HS65_LH_AO222X4 U8754 ( .A(n7896), .B(\u_DataPath/pc_4_i [25]), .C(n7893), 
        .D(n9415), .E(n9199), .F(n7887), .Z(n8647) );
  HS65_LH_AO222X4 U8755 ( .A(n7895), .B(\u_DataPath/pc_4_i [15]), .C(n7892), 
        .D(n9418), .E(n8930), .F(n7888), .Z(n8657) );
  HS65_LH_AO222X4 U8756 ( .A(n7895), .B(\u_DataPath/pc_4_i [13]), .C(n7892), 
        .D(n9413), .E(n8919), .F(n7888), .Z(n8659) );
  HS65_LH_AO222X4 U8757 ( .A(n7895), .B(\u_DataPath/pc_4_i [20]), .C(n7892), 
        .D(n9404), .E(n8926), .F(n7887), .Z(n8652) );
  HS65_LH_NAND2X2 U8758 ( .A(n2733), .B(\u_DataPath/cw_memwb_i [2]), .Z(n8061)
         );
  HS65_LH_NOR2X2 U8759 ( .A(n8107), .B(rst), .Z(
        \u_DataPath/regfile_addr_out_towb_i [4]) );
  HS65_LH_CNIVX3 U8760 ( .A(n8763), .Z(n8108) );
  HS65_LH_AO22X4 U8761 ( .A(n9267), .B(n8067), .C(n8967), .D(n8066), .Z(
        \u_DataPath/RFaddr_out_memwb_i [2]) );
  HS65_LH_AO22X4 U8762 ( .A(n9183), .B(n8067), .C(n8942), .D(n8066), .Z(
        \u_DataPath/RFaddr_out_memwb_i [0]) );
  HS65_LH_AO22X4 U8763 ( .A(n9145), .B(n8067), .C(n8968), .D(n8066), .Z(
        \u_DataPath/RFaddr_out_memwb_i [4]) );
  HS65_LH_AO22X4 U8764 ( .A(n9181), .B(n8067), .C(n9077), .D(n8066), .Z(
        \u_DataPath/RFaddr_out_memwb_i [3]) );
  HS65_LH_AOI22X1 U8765 ( .A(n8868), .B(n9184), .C(n9365), .D(n9057), .Z(n8416) );
  HS65_LH_NAND3X2 U8766 ( .A(n2733), .B(n8715), .C(\u_DataPath/cw_to_ex_i [15]), .Z(n8428) );
  HS65_LH_AOI22X1 U8768 ( .A(n8868), .B(n9170), .C(n9365), .D(n9020), .Z(n8317) );
  HS65_LH_CNIVX3 U8769 ( .A(n9207), .Z(n7119) );
  HS65_LH_AOI22X1 U8770 ( .A(n8868), .B(n9172), .C(n9369), .D(n8987), .Z(n8328) );
  HS65_LH_OAI21X3 U8771 ( .A(n9189), .B(n8902), .C(n8375), .Z(
        \u_DataPath/dataOut_exe_i [27]) );
  HS65_LH_AOI22X1 U8772 ( .A(n8868), .B(n9182), .C(n9366), .D(n8996), .Z(n8375) );
  HS65_LL_OAI21X12 U8773 ( .A(n3009), .B(n8140), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N140 ) );
  HS65_LL_OAI21X12 U8774 ( .A(n8140), .B(n2773), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N141 ) );
  HS65_LL_OAI21X12 U8775 ( .A(n8140), .B(n8147), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N143 ) );
  HS65_LL_OAI21X12 U8776 ( .A(n8140), .B(n3010), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N145 ) );
  HS65_LHS_XOR2X3 U8777 ( .A(n6037), .B(n6089), .Z(
        \u_DataPath/u_execute/resAdd1_i [6]) );
  HS65_LHS_XOR2X3 U8778 ( .A(n6012), .B(n6065), .Z(
        \u_DataPath/u_execute/resAdd1_i [18]) );
  HS65_LHS_XOR2X3 U8779 ( .A(n6025), .B(n6024), .Z(
        \u_DataPath/u_execute/resAdd1_i [17]) );
  HS65_LHS_XOR2X3 U8780 ( .A(n6004), .B(n6003), .Z(
        \u_DataPath/u_execute/resAdd1_i [20]) );
  HS65_LH_NAND3AX3 U8781 ( .A(n5693), .B(n5692), .C(n5691), .Z(n8503) );
  HS65_LHS_XOR2X3 U8782 ( .A(n6032), .B(n6077), .Z(
        \u_DataPath/u_execute/resAdd1_i [8]) );
  HS65_LH_NAND2X2 U8783 ( .A(n6110), .B(n6109), .Z(n6112) );
  HS65_LH_NAND2X2 U8784 ( .A(n6106), .B(n6105), .Z(n6108) );
  HS65_LHS_XOR2X3 U8786 ( .A(n6044), .B(n6043), .Z(
        \u_DataPath/u_execute/resAdd1_i [5]) );
  HS65_LHS_XOR2X3 U8787 ( .A(n6018), .B(n6017), .Z(
        \u_DataPath/u_execute/resAdd1_i [21]) );
  HS65_LHS_XOR2X3 U8788 ( .A(n5994), .B(n5993), .Z(
        \u_DataPath/u_execute/resAdd1_i [13]) );
  HS65_LH_CNIVX3 U8789 ( .A(n6125), .Z(n8513) );
  HS65_LH_AO22X9 U8790 ( .A(n9258), .B(n9188), .C(n9133), .D(n8999), .Z(
        \u_DataPath/jump_address_i [30]) );
  HS65_LHS_XNOR2X3 U8791 ( .A(n6072), .B(n6071), .Z(
        \u_DataPath/u_execute/resAdd1_i [10]) );
  HS65_LH_AOI21X2 U8792 ( .A(n2866), .B(n8537), .C(n8536), .Z(
        \u_DataPath/mem_writedata_out_i [19]) );
  HS65_LHS_XOR2X3 U8793 ( .A(n5986), .B(n5985), .Z(
        \u_DataPath/u_execute/resAdd1_i [11]) );
  HS65_LH_NOR4ABX2 U8794 ( .A(n6224), .B(n6223), .C(n6222), .D(n6221), .Z(
        n8377) );
  HS65_LHS_XOR2X3 U8795 ( .A(n5970), .B(n5969), .Z(
        \u_DataPath/u_execute/resAdd1_i [15]) );
  HS65_LHS_XNOR2X3 U8796 ( .A(n6060), .B(n6059), .Z(
        \u_DataPath/u_execute/resAdd1_i [14]) );
  HS65_LH_NOR4ABX2 U8797 ( .A(n6393), .B(n6392), .C(n6391), .D(n6390), .Z(
        n8309) );
  HS65_LH_NOR4ABX2 U8798 ( .A(n6264), .B(n6263), .C(n6262), .D(n6261), .Z(
        n8347) );
  HS65_LH_NOR4ABX2 U8799 ( .A(n6534), .B(n6533), .C(n6532), .D(n6531), .Z(
        n8325) );
  HS65_LH_NOR4ABX2 U8801 ( .A(n6594), .B(n6593), .C(n6592), .D(n6591), .Z(
        n8174) );
  HS65_LH_NOR4ABX2 U8802 ( .A(n6413), .B(n6412), .C(n6411), .D(n6410), .Z(
        n8296) );
  HS65_LH_CNIVX3 U8803 ( .A(n9214), .Z(n7727) );
  HS65_LH_NOR4ABX2 U8804 ( .A(n6514), .B(n6513), .C(n6512), .D(n6511), .Z(
        n8320) );
  HS65_LH_NOR4ABX2 U8805 ( .A(n6244), .B(n6243), .C(n6242), .D(n6241), .Z(
        n8361) );
  HS65_LH_AOI22X1 U8806 ( .A(n8868), .B(n9174), .C(n9368), .D(n8975), .Z(n8359) );
  HS65_LH_NOR4ABX2 U8807 ( .A(n6554), .B(n6553), .C(n6552), .D(n6551), .Z(
        n8292) );
  HS65_LH_NOR4ABX2 U8808 ( .A(n6454), .B(n6453), .C(n6452), .D(n6451), .Z(
        n8303) );
  HS65_LH_CNIVX3 U8809 ( .A(n9227), .Z(n7709) );
  HS65_LH_CNIVX3 U8810 ( .A(n9228), .Z(n7732) );
  HS65_LH_NOR4ABX2 U8811 ( .A(n6950), .B(n6949), .C(n6948), .D(n6947), .Z(
        n8414) );
  HS65_LH_AOI22X1 U8813 ( .A(n8868), .B(n9176), .C(n9369), .D(n8983), .Z(n8369) );
  HS65_LH_CNIVX3 U8814 ( .A(n9209), .Z(n7121) );
  HS65_LH_NOR4ABX2 U8815 ( .A(n6926), .B(n6925), .C(n6924), .D(n6923), .Z(
        n8418) );
  HS65_LH_AOI22X1 U8816 ( .A(n8868), .B(n9178), .C(n9365), .D(n8938), .Z(n7856) );
  HS65_LH_CBI4I1X3 U8817 ( .A(n2874), .B(n8724), .C(n7846), .D(n8566), .Z(
        n8493) );
  HS65_LH_AO22X9 U8818 ( .A(n8872), .B(n9188), .C(n9133), .D(n9041), .Z(
        \u_DataPath/jump_address_i [4]) );
  HS65_LH_NOR4ABX2 U8819 ( .A(n6649), .B(n6648), .C(n6647), .D(n6646), .Z(
        n8430) );
  HS65_LH_CNIVX3 U8820 ( .A(n9219), .Z(n7726) );
  HS65_LH_NOR4ABX2 U8821 ( .A(n6474), .B(n6473), .C(n6472), .D(n6471), .Z(
        n8274) );
  HS65_LHS_XNOR2X3 U8822 ( .A(n7719), .B(n7781), .Z(
        \u_DataPath/u_execute/link_value_i [8]) );
  HS65_LH_CNIVX3 U8823 ( .A(n9229), .Z(n7719) );
  HS65_LH_NOR4ABX2 U8824 ( .A(n6866), .B(n6865), .C(n6864), .D(n6863), .Z(
        n8411) );
  HS65_LH_AOI22X1 U8825 ( .A(n8868), .B(n8912), .C(n9366), .D(n9046), .Z(n8409) );
  HS65_LH_NOR4ABX2 U8826 ( .A(n6184), .B(n6183), .C(n6182), .D(n6181), .Z(
        n8357) );
  HS65_LHS_XOR2X3 U8828 ( .A(n7715), .B(n7714), .Z(n5690) );
  HS65_LH_NOR4ABX2 U8829 ( .A(n6906), .B(n6905), .C(n6904), .D(n6903), .Z(
        n8407) );
  HS65_LH_AOI22X1 U8830 ( .A(n8868), .B(n9036), .C(n9366), .D(n9017), .Z(n8405) );
  HS65_LH_AOI21X2 U8831 ( .A(n2874), .B(n8490), .C(n8489), .Z(
        \u_DataPath/mem_writedata_out_i [2]) );
  HS65_LH_AO22X9 U8832 ( .A(n9188), .B(n9021), .C(n9133), .D(n8945), .Z(
        \u_DataPath/jump_address_i [2]) );
  HS65_LHS_XOR2X3 U8833 ( .A(n6052), .B(n6101), .Z(
        \u_DataPath/u_execute/resAdd1_i [2]) );
  HS65_LH_NOR4ABX2 U8834 ( .A(n6574), .B(n6573), .C(n6572), .D(n6571), .Z(
        n8173) );
  HS65_LH_NOR4ABX2 U8835 ( .A(n6669), .B(n6668), .C(n6667), .D(n6666), .Z(
        n8455) );
  HS65_LH_MX41X4 U8836 ( .D0(n8441), .S0(n9280), .D1(n8440), .S1(n9295), .D2(
        n9302), .S2(n8439), .D3(n8438), .S3(n9287), .Z(
        \u_DataPath/from_mem_data_out_i [6]) );
  HS65_LH_MX41X4 U8837 ( .D0(n8441), .S0(n9279), .D1(n8440), .S1(n9294), .D2(
        n9301), .S2(n8439), .D3(n8438), .S3(n9286), .Z(
        \u_DataPath/from_mem_data_out_i [5]) );
  HS65_LH_MX41X4 U8838 ( .D0(n8441), .S0(n9278), .D1(n8440), .S1(n9293), .D2(
        n9300), .S2(n8439), .D3(n8438), .S3(n9285), .Z(
        \u_DataPath/from_mem_data_out_i [4]) );
  HS65_LH_MX41X4 U8839 ( .D0(n8441), .S0(n9277), .D1(n8440), .S1(n9292), .D2(
        n9299), .S2(n8439), .D3(n8438), .S3(n9284), .Z(
        \u_DataPath/from_mem_data_out_i [3]) );
  HS65_LH_MX41X4 U8840 ( .D0(n8441), .S0(n9276), .D1(n8440), .S1(n9291), .D2(
        n9298), .S2(n8439), .D3(n8438), .S3(n9283), .Z(
        \u_DataPath/from_mem_data_out_i [2]) );
  HS65_LH_AO22X9 U8841 ( .A(n9133), .B(n8935), .C(n9188), .D(n9105), .Z(
        \u_DataPath/jump_address_i [1]) );
  HS65_LH_NOR4ABX2 U8843 ( .A(n6616), .B(n6615), .C(n6614), .D(n6613), .Z(
        n8167) );
  HS65_LH_OR2X4 U8846 ( .A(n9035), .B(n9115), .Z(n5918) );
  HS65_LH_NOR4ABX2 U8847 ( .A(n6434), .B(n6433), .C(n6432), .D(n6431), .Z(
        n8169) );
  HS65_LH_NOR4ABX2 U8848 ( .A(n6886), .B(n6885), .C(n6884), .D(n6883), .Z(
        n8421) );
  HS65_LH_AO22X4 U8849 ( .A(n8757), .B(n9138), .C(n9320), .D(n9153), .Z(
        \u_DataPath/jaddr_i [17]) );
  HS65_LH_NOR2X2 U8850 ( .A(n8164), .B(rst), .Z(\u_DataPath/rs_ex_i [1]) );
  HS65_LH_NOR2X2 U8851 ( .A(n8165), .B(rst), .Z(\u_DataPath/rs_ex_i [2]) );
  HS65_LH_AO22X4 U8852 ( .A(n8756), .B(n9252), .C(n9328), .D(n9153), .Z(
        \u_DataPath/jaddr_i [25]) );
  HS65_LH_NAND2AX4 U8853 ( .A(n8480), .B(\u_DataPath/u_idexreg/N10 ), .Z(n8136) );
  HS65_LH_NAND2AX4 U8854 ( .A(n8480), .B(\u_DataPath/u_idexreg/N16 ), .Z(n8111) );
  HS65_LH_NAND2AX4 U8855 ( .A(n8480), .B(\u_DataPath/cw_exmem_i [5]), .Z(n8113) );
  HS65_LH_NAND2AX4 U8856 ( .A(n8480), .B(\u_DataPath/u_idexreg/N15 ), .Z(n8112) );
  HS65_LH_NAND2AX4 U8857 ( .A(n8480), .B(\u_DataPath/cw_exmem_i [4]), .Z(n8109) );
  HS65_LH_NOR4ABX4 U8858 ( .A(opcode_i[1]), .B(n8116), .C(n8056), .D(n8117), 
        .Z(\u_DataPath/cw_to_ex_i [17]) );
  HS65_LH_NAND2AX4 U8859 ( .A(n8480), .B(\u_DataPath/cw_exmem_i [6]), .Z(n8110) );
  HS65_LH_NAND2AX4 U8860 ( .A(n8480), .B(n9052), .Z(n8481) );
  HS65_LH_NAND2AX4 U8861 ( .A(n8480), .B(n9048), .Z(n8233) );
  HS65_LH_NOR2X2 U8862 ( .A(n8152), .B(rst), .Z(\u_DataPath/idex_rt_i [0]) );
  HS65_LH_AO22X4 U8863 ( .A(n8754), .B(n9138), .C(n9319), .D(n9153), .Z(
        \u_DataPath/jaddr_i [16]) );
  HS65_LH_AND2X4 U8864 ( .A(n2733), .B(\u_DataPath/toPC2_i [28]), .Z(
        \u_DataPath/branch_target_i [28]) );
  HS65_LH_CNIVX3 U8865 ( .A(n5743), .Z(n5744) );
  HS65_LH_AND2X4 U8866 ( .A(n2733), .B(\u_DataPath/toPC2_i [26]), .Z(
        \u_DataPath/branch_target_i [26]) );
  HS65_LHS_XOR2X3 U8867 ( .A(n5810), .B(n5809), .Z(\u_DataPath/toPC2_i [20])
         );
  HS65_LHS_XOR2X3 U8868 ( .A(n5804), .B(n5803), .Z(\u_DataPath/toPC2_i [19])
         );
  HS65_LHS_XOR2X3 U8869 ( .A(n5816), .B(n5815), .Z(\u_DataPath/toPC2_i [18])
         );
  HS65_LHS_XOR2X3 U8870 ( .A(n5823), .B(n5822), .Z(\u_DataPath/toPC2_i [17])
         );
  HS65_LHS_XOR2X3 U8871 ( .A(n5766), .B(n5765), .Z(\u_DataPath/toPC2_i [15])
         );
  HS65_LH_AOI12X2 U8872 ( .A(n6057), .B(n5864), .C(n5764), .Z(n5765) );
  HS65_LHS_XNOR2X3 U8873 ( .A(n5865), .B(n5864), .Z(\u_DataPath/toPC2_i [14])
         );
  HS65_LHS_XOR2X3 U8874 ( .A(n5794), .B(n5793), .Z(\u_DataPath/toPC2_i [13])
         );
  HS65_LHS_XOR2X3 U8875 ( .A(n5785), .B(n5784), .Z(\u_DataPath/toPC2_i [11])
         );
  HS65_LHS_XNOR2X3 U8876 ( .A(n5873), .B(n5872), .Z(\u_DataPath/toPC2_i [10])
         );
  HS65_LHS_XOR2X3 U8877 ( .A(n5830), .B(n5878), .Z(\u_DataPath/toPC2_i [8]) );
  HS65_LHS_XOR2X3 U8879 ( .A(n5835), .B(n5886), .Z(\u_DataPath/toPC2_i [6]) );
  HS65_LHS_XOR2X3 U8881 ( .A(n5842), .B(n5841), .Z(\u_DataPath/toPC2_i [5]) );
  HS65_LHS_XOR2X3 U8882 ( .A(n5845), .B(n5898), .Z(\u_DataPath/toPC2_i [2]) );
  HS65_LL_NOR4ABX2 U8885 ( .A(n7243), .B(n7242), .C(n7241), .D(n7240), .Z(
        n8178) );
  HS65_LL_NOR4ABX2 U8887 ( .A(n7342), .B(n7341), .C(n7340), .D(n7339), .Z(
        n8315) );
  HS65_LL_NOR4ABX2 U8889 ( .A(n7263), .B(n7262), .C(n7261), .D(n7260), .Z(
        n8310) );
  HS65_LLS_XNOR2X3 U8892 ( .A(n4422), .B(n4421), .Z(n4423) );
  HS65_LL_AND2X4 U8893 ( .A(n4714), .B(n8515), .Z(n3261) );
  HS65_LH_AOI22X1 U8894 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][4] ), .B(n6754), 
        .C(n6684), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][4] ), .Z(n7355)
         );
  HS65_LH_NOR2X6 U8895 ( .A(n6353), .B(n6332), .Z(n2889) );
  HS65_LH_NOR2X6 U8896 ( .A(n6350), .B(n6332), .Z(n2890) );
  HS65_LH_NOR2X6 U8897 ( .A(n6349), .B(n2878), .Z(n2891) );
  HS65_LH_AOI22X1 U8898 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][23] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ), .D(
        n6171), .Z(n6234) );
  HS65_LH_AOI22X1 U8899 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][27] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][27] ), .D(
        n6171), .Z(n6214) );
  HS65_LL_NOR3AX9 U8901 ( .A(n3344), .B(n3343), .C(n3342), .Z(\lte_x_59/B[4] )
         );
  HS65_LH_NOR2X2 U8902 ( .A(n3474), .B(n3359), .Z(n5298) );
  HS65_LL_NAND4ABX3 U8903 ( .A(n3824), .B(n3823), .C(n3822), .D(n3821), .Z(
        n4840) );
  HS65_LH_NOR2X2 U8904 ( .A(\lte_x_59/B[24] ), .B(n3382), .Z(n5426) );
  HS65_LH_AND3X4 U8905 ( .A(n4836), .B(\sub_x_53/A[2] ), .C(n4552), .Z(n2901)
         );
  HS65_LL_NOR2AX3 U8906 ( .A(n3554), .B(n3553), .Z(n3555) );
  HS65_LL_AND2X4 U8907 ( .A(n9205), .B(n7307), .Z(n2908) );
  HS65_LL_AND2X4 U8908 ( .A(n2963), .B(n2962), .Z(n2912) );
  HS65_LL_OR2X4 U8909 ( .A(n8798), .B(n3403), .Z(n2913) );
  HS65_LL_AND2X4 U8910 ( .A(n4289), .B(n4211), .Z(n2914) );
  HS65_LL_AND2X4 U8911 ( .A(n4714), .B(n8530), .Z(n2919) );
  HS65_LL_AND2X4 U8912 ( .A(n3327), .B(n9145), .Z(n2922) );
  HS65_LH_AND2X4 U8913 ( .A(n4717), .B(n9181), .Z(n2923) );
  HS65_LH_IVX9 U8915 ( .A(n7802), .Z(n8390) );
  HS65_LLS_XNOR2X3 U8916 ( .A(n3008), .B(n8942), .Z(n2953) );
  HS65_LLS_XNOR2X3 U8917 ( .A(n7086), .B(n2950), .Z(n2951) );
  HS65_LL_AND2ABX18 U8919 ( .A(n7638), .B(n2974), .Z(write_byte) );
  HS65_LL_AND2X18 U8920 ( .A(n8879), .B(write_op), .Z(Data_in[4]) );
  HS65_LL_NOR2AX25 U8921 ( .A(\u_DataPath/dataOut_exe_i [31]), .B(n3116), .Z(
        Address_toRAM[29]) );
  HS65_LL_NOR2AX25 U8922 ( .A(\u_DataPath/dataOut_exe_i [9]), .B(n2986), .Z(
        Address_toRAM[7]) );
  HS65_LL_NOR2AX25 U8923 ( .A(\u_DataPath/dataOut_exe_i [7]), .B(n2986), .Z(
        Address_toRAM[5]) );
  HS65_LL_NOR2AX25 U8924 ( .A(\u_DataPath/dataOut_exe_i [14]), .B(n2986), .Z(
        Address_toRAM[12]) );
  HS65_LL_NOR2AX25 U8925 ( .A(\u_DataPath/dataOut_exe_i [16]), .B(n2986), .Z(
        Address_toRAM[14]) );
  HS65_LL_NOR2AX25 U8926 ( .A(n8738), .B(n2994), .Z(Data_in[16]) );
  HS65_LL_NOR2AX25 U8927 ( .A(n8739), .B(n2994), .Z(Data_in[14]) );
  HS65_LL_NOR2AX25 U8928 ( .A(n8730), .B(n2994), .Z(Data_in[12]) );
  HS65_LL_NOR2AX25 U8929 ( .A(n8735), .B(n2994), .Z(Data_in[11]) );
  HS65_LL_NOR2AX25 U8930 ( .A(n8741), .B(n2994), .Z(Data_in[10]) );
  HS65_LL_NOR2AX25 U8931 ( .A(n8734), .B(n2994), .Z(Data_in[15]) );
  HS65_LL_NOR2AX25 U8932 ( .A(n8740), .B(n2994), .Z(Data_in[17]) );
  HS65_LL_NOR2AX25 U8933 ( .A(n8746), .B(n2994), .Z(Data_in[21]) );
  HS65_LL_NOR2AX25 U8934 ( .A(n8747), .B(n2994), .Z(Data_in[20]) );
  HS65_LL_NOR2AX25 U8935 ( .A(\u_DataPath/dataOut_exe_i [15]), .B(n2986), .Z(
        Address_toRAM[13]) );
  HS65_LL_NOR2AX25 U8936 ( .A(\u_DataPath/dataOut_exe_i [17]), .B(n2986), .Z(
        Address_toRAM[15]) );
  HS65_LL_NOR2AX25 U8937 ( .A(\u_DataPath/dataOut_exe_i [26]), .B(n3116), .Z(
        Address_toRAM[24]) );
  HS65_LH_IVX2 U8939 ( .A(n7086), .Z(n3011) );
  HS65_LL_AND2X18 U8940 ( .A(n9018), .B(write_op), .Z(Data_in[0]) );
  HS65_LH_OAI22X1 U8941 ( .A(n3285), .B(n4712), .C(n3288), .D(n9401), .Z(n8484) );
  HS65_LH_MUXI21X2 U8942 ( .D0(n3018), .D1(n9379), .S0(n3404), .Z(n8243) );
  HS65_LH_MUXI21X2 U8943 ( .D0(n3020), .D1(n9393), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8374) );
  HS65_LH_NAND2X7 U8944 ( .A(\u_DataPath/cw_memwb_i [2]), .B(n3035), .Z(n3044)
         );
  HS65_LLS_XNOR2X3 U8945 ( .A(n8762), .B(n8911), .Z(n3038) );
  HS65_LH_MUXI21X2 U8946 ( .D0(n3047), .D1(n9392), .S0(n3404), .Z(n8380) );
  HS65_LH_AND2X4 U8947 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n3407), .Z(
        n3068) );
  HS65_LH_NOR2X6 U8948 ( .A(n8831), .B(n3341), .Z(n3073) );
  HS65_LH_NOR2X6 U8949 ( .A(n8826), .B(n3341), .Z(n3076) );
  HS65_LH_MUXI21X2 U8950 ( .D0(n3079), .D1(n9398), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8332) );
  HS65_LH_MUXI21X2 U8951 ( .D0(n3084), .D1(n9391), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8387) );
  HS65_LH_NOR2X6 U8952 ( .A(n8851), .B(n3341), .Z(n3091) );
  HS65_LH_MUXI21X2 U8953 ( .D0(n3088), .D1(n9382), .S0(n3404), .Z(n8389) );
  HS65_LH_MUXI21X2 U8954 ( .D0(n3093), .D1(n9390), .S0(n3404), .Z(n8355) );
  HS65_LH_NOR2X6 U8955 ( .A(n8855), .B(n3403), .Z(n3106) );
  HS65_LH_MUXI21X2 U8956 ( .D0(n3103), .D1(n9378), .S0(n3404), .Z(n8266) );
  HS65_LL_AO112X18 U8957 ( .A(n8578), .B(n3112), .C(n2879), .D(n8577), .Z(
        read_op) );
  HS65_LL_OR2ABX18 U8958 ( .A(n8576), .B(n8575), .Z(nibble[1]) );
  HS65_LL_NOR2AX25 U8959 ( .A(\u_DataPath/dataOut_exe_i [6]), .B(n2986), .Z(
        Address_toRAM[4]) );
  HS65_LL_NOR2AX25 U8960 ( .A(\u_DataPath/dataOut_exe_i [5]), .B(n2986), .Z(
        Address_toRAM[3]) );
  HS65_LL_NOR2AX25 U8961 ( .A(\u_DataPath/dataOut_exe_i [3]), .B(n2986), .Z(
        Address_toRAM[1]) );
  HS65_LL_NOR2AX25 U8962 ( .A(\u_DataPath/dataOut_exe_i [19]), .B(n3116), .Z(
        Address_toRAM[17]) );
  HS65_LL_NOR2AX25 U8963 ( .A(\u_DataPath/dataOut_exe_i [18]), .B(n3116), .Z(
        Address_toRAM[16]) );
  HS65_LL_NOR2AX25 U8964 ( .A(\u_DataPath/dataOut_exe_i [2]), .B(n3116), .Z(
        Address_toRAM[0]) );
  HS65_LL_NOR2AX25 U8965 ( .A(n8733), .B(n3115), .Z(Data_in[26]) );
  HS65_LL_NOR2AX25 U8966 ( .A(n9085), .B(n3115), .Z(Data_in[25]) );
  HS65_LL_NOR2AX25 U8967 ( .A(n8732), .B(n3115), .Z(Data_in[24]) );
  HS65_LL_AND2ABX18 U8968 ( .A(n8574), .B(n3116), .Z(Address_toRAM[2]) );
  HS65_LH_IVX40 U8969 ( .A(n3126), .Z(addr_to_iram[1]) );
  HS65_LL_AND2X18 U8970 ( .A(n8731), .B(write_op), .Z(Data_in[5]) );
  HS65_LL_AND2X18 U8971 ( .A(n8744), .B(write_op), .Z(Data_in[1]) );
  HS65_LL_AND2X18 U8972 ( .A(n8745), .B(write_op), .Z(Data_in[7]) );
  HS65_LL_AND2X18 U8973 ( .A(n8725), .B(write_op), .Z(Data_in[3]) );
  HS65_LL_AND2X18 U8974 ( .A(n8873), .B(write_op), .Z(Data_in[2]) );
  HS65_LL_AND2X18 U8975 ( .A(n8743), .B(write_op), .Z(Data_in[6]) );
  HS65_LH_BFX18 U8978 ( .A(n9376), .Z(n4714) );
  HS65_LH_NOR2X6 U8980 ( .A(n3572), .B(n3575), .Z(n3751) );
  HS65_LH_MUXI21X2 U8981 ( .D0(n7877), .D1(n9388), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8316) );
  HS65_LL_MUXI21X2 U8982 ( .D0(n3185), .D1(n9387), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8323) );
  HS65_LH_IVX9 U8983 ( .A(n5005), .Z(n3371) );
  HS65_LH_NOR2X6 U8984 ( .A(n8822), .B(n3403), .Z(n3200) );
  HS65_LH_NOR2X6 U8985 ( .A(\sub_x_53/A[17] ), .B(n2870), .Z(n3515) );
  HS65_LH_NOR2X6 U8986 ( .A(n8860), .B(n3403), .Z(n3214) );
  HS65_LH_NOR2X2 U8987 ( .A(n8265), .B(n8262), .Z(n3219) );
  HS65_LH_MUXI21X2 U8989 ( .D0(n3248), .D1(n9397), .S0(n3404), .Z(n8339) );
  HS65_LH_MUXI21X2 U8990 ( .D0(n3259), .D1(n9381), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8255) );
  HS65_LH_MUXI21X2 U8991 ( .D0(n8909), .D1(
        \u_DataPath/from_mem_data_out_i [15]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n8306) );
  HS65_LH_NOR2X6 U8992 ( .A(n8840), .B(n3290), .Z(n3292) );
  HS65_LL_OAI22X3 U8993 ( .A(n3333), .B(\u_DataPath/dataOut_exe_i [2]), .C(
        n8488), .D(n3340), .Z(n3295) );
  HS65_LH_NAND2X7 U8994 ( .A(n3296), .B(n7802), .Z(n8487) );
  HS65_LH_AND2X4 U8995 ( .A(n3309), .B(n3308), .Z(n3311) );
  HS65_LH_NOR2X6 U8996 ( .A(n8857), .B(n3403), .Z(n3320) );
  HS65_LH_AND2X4 U8998 ( .A(n2896), .B(n3337), .Z(n7863) );
  HS65_LH_NAND2X7 U8999 ( .A(\lte_x_59/B[18] ), .B(n3371), .Z(n5272) );
  HS65_LH_NAND2X7 U9000 ( .A(n2849), .B(n3372), .Z(n5270) );
  HS65_LH_MUX21I1X3 U9001 ( .D0(n3402), .D1(n5183), .S0(n5088), .Z(n4457) );
  HS65_LH_NOR2X6 U9002 ( .A(n8823), .B(n3403), .Z(n3411) );
  HS65_LL_NOR2AX3 U9003 ( .A(n2866), .B(n3418), .Z(n7846) );
  HS65_LH_AOI22X1 U9004 ( .A(\sub_x_53/A[23] ), .B(n4587), .C(n2864), .D(
        \lte_x_59/B[21] ), .Z(n3435) );
  HS65_LH_NOR2X2 U9005 ( .A(n4726), .B(n2893), .Z(n3439) );
  HS65_LH_NAND3X2 U9006 ( .A(n4551), .B(n4836), .C(n4949), .Z(n3444) );
  HS65_LH_AOI22X1 U9007 ( .A(\sub_x_53/A[27] ), .B(n4587), .C(n3789), .D(
        \sub_x_53/A[25] ), .Z(n3445) );
  HS65_LH_NAND2X7 U9008 ( .A(n5321), .B(n5088), .Z(n4838) );
  HS65_LH_OAI21X3 U9009 ( .A(n3272), .B(n2857), .C(n3839), .Z(n3459) );
  HS65_LH_NOR2AX3 U9010 ( .A(n3469), .B(n3468), .Z(n3512) );
  HS65_LH_CNIVX3 U9012 ( .A(n3617), .Z(n3494) );
  HS65_LH_NAND2X2 U9014 ( .A(\lte_x_59/B[9] ), .B(n4551), .Z(n3526) );
  HS65_LH_NAND3X2 U9015 ( .A(\sub_x_53/A[17] ), .B(n3582), .C(n5001), .Z(n3531) );
  HS65_LH_CBI4I1X3 U9016 ( .A(n9352), .B(n5001), .C(\sub_x_53/A[17] ), .D(
        n5647), .Z(n3530) );
  HS65_LH_OAI21X3 U9017 ( .A(n5621), .B(n4889), .C(n3604), .Z(n3605) );
  HS65_LH_NOR2AX3 U9018 ( .A(\sub_x_53/A[2] ), .B(n2857), .Z(n3641) );
  HS65_LH_OA12X9 U9019 ( .A(n5129), .B(n4811), .C(n4794), .Z(n3642) );
  HS65_LH_NOR2X6 U9020 ( .A(n2840), .B(n3756), .Z(n4507) );
  HS65_LH_NAND3X2 U9022 ( .A(n4836), .B(n5624), .C(n4504), .Z(n3653) );
  HS65_LH_AOI22X1 U9023 ( .A(n2849), .B(n4588), .C(n4587), .D(\lte_x_59/B[18] ), .Z(n3663) );
  HS65_LH_AOI21X2 U9024 ( .A(n5618), .B(n5228), .C(n3668), .Z(n3677) );
  HS65_LL_NOR3X1 U9025 ( .A(n3681), .B(n3680), .C(n3679), .Z(n3695) );
  HS65_LLS_XNOR2X3 U9026 ( .A(n3692), .B(n3691), .Z(n3693) );
  HS65_LLS_XNOR2X3 U9027 ( .A(n3708), .B(n3707), .Z(n3746) );
  HS65_LH_OAI21X3 U9028 ( .A(n5240), .B(n4855), .C(n3714), .Z(n3715) );
  HS65_LH_CNIVX3 U9029 ( .A(n5608), .Z(n3734) );
  HS65_LLS_XNOR2X3 U9030 ( .A(n3755), .B(n3754), .Z(n3813) );
  HS65_LH_MUXI21X2 U9031 ( .D0(n4726), .D1(n2840), .S0(n3756), .Z(n4491) );
  HS65_LHS_XNOR2X3 U9032 ( .A(n2853), .B(n5567), .Z(n4751) );
  HS65_LH_OAI21X3 U9033 ( .A(n4986), .B(n3756), .C(n3768), .Z(n3769) );
  HS65_LH_NAND3X2 U9034 ( .A(n3582), .B(n2853), .C(n5567), .Z(n3776) );
  HS65_LH_NAND2X2 U9035 ( .A(n5647), .B(n2853), .Z(n3775) );
  HS65_LH_AND2X4 U9036 ( .A(\lte_x_59/B[7] ), .B(n3789), .Z(n4465) );
  HS65_LH_NAND2X2 U9037 ( .A(n5207), .B(n5660), .Z(n3791) );
  HS65_LH_CBI4I1X3 U9038 ( .A(n3582), .B(n5048), .C(n5647), .D(n3521), .Z(
        n3825) );
  HS65_LH_NAND2X7 U9039 ( .A(n4836), .B(n4550), .Z(n5201) );
  HS65_LHS_XNOR2X6 U9041 ( .A(n3848), .B(n3847), .Z(n3849) );
  HS65_LH_CNIVX3 U9042 ( .A(n5143), .Z(n3874) );
  HS65_LH_NAND3X2 U9043 ( .A(n4512), .B(n3426), .C(n3872), .Z(n3873) );
  HS65_LH_NAND3X2 U9044 ( .A(n4949), .B(n3426), .C(n4176), .Z(n3922) );
  HS65_LH_CNIVX3 U9045 ( .A(n4754), .Z(n3975) );
  HS65_LH_NAND3X2 U9046 ( .A(n4192), .B(n5032), .C(n3969), .Z(n3972) );
  HS65_LH_NAND2X2 U9047 ( .A(n9352), .B(n5104), .Z(n3971) );
  HS65_LH_IVX9 U9048 ( .A(n4287), .Z(n7729) );
  HS65_LH_AND2X4 U9049 ( .A(n4041), .B(n4037), .Z(n4043) );
  HS65_LHS_XNOR2X3 U9050 ( .A(n4674), .B(n2842), .Z(n4740) );
  HS65_LH_AOI22X1 U9051 ( .A(n4516), .B(n5239), .C(n4508), .D(n4614), .Z(n4179) );
  HS65_LH_NAND2X2 U9052 ( .A(n3426), .B(n4176), .Z(n4178) );
  HS65_LH_AOI22X1 U9053 ( .A(\sub_x_53/A[30] ), .B(n4587), .C(n4351), .D(
        \sub_x_53/A[29] ), .Z(n4182) );
  HS65_LH_CNIVX3 U9054 ( .A(n4738), .Z(n4199) );
  HS65_LLS_XNOR2X3 U9055 ( .A(n5005), .B(\lte_x_59/B[18] ), .Z(n4744) );
  HS65_LH_CBI4I1X3 U9056 ( .A(n5648), .B(n5005), .C(n5647), .D(
        \lte_x_59/B[18] ), .Z(n4270) );
  HS65_LL_AOI22X1 U9057 ( .A(n8868), .B(n9038), .C(n9366), .D(n8972), .Z(n7843) );
  HS65_LLS_XNOR2X3 U9058 ( .A(n4339), .B(n4338), .Z(n4367) );
  HS65_LH_NAND2X2 U9059 ( .A(n4340), .B(n4341), .Z(n4343) );
  HS65_LH_OAI22X1 U9060 ( .A(n2854), .B(n4795), .C(n2857), .D(n4724), .Z(n4350) );
  HS65_LHS_XNOR2X3 U9061 ( .A(\lte_x_59/B[21] ), .B(n5418), .Z(n4737) );
  HS65_LH_NAND2X2 U9062 ( .A(n5207), .B(n4872), .Z(n4392) );
  HS65_LH_CBI4I1X3 U9063 ( .A(n5648), .B(n5418), .C(n5647), .D(
        \lte_x_59/B[21] ), .Z(n4396) );
  HS65_LL_NAND3X2 U9064 ( .A(n4400), .B(n4399), .C(n4398), .Z(n4401) );
  HS65_LHS_XNOR2X3 U9065 ( .A(\lte_x_59/B[4] ), .B(n5032), .Z(n4749) );
  HS65_LH_CBI4I1X3 U9066 ( .A(n5648), .B(n2872), .C(n3443), .D(\lte_x_59/B[4] ), .Z(n4459) );
  HS65_LH_NOR2X2 U9067 ( .A(n4513), .B(n4838), .Z(n4514) );
  HS65_LH_OAI22X1 U9068 ( .A(n4725), .B(n4583), .C(n5129), .D(n4724), .Z(n4523) );
  HS65_LHS_XNOR2X6 U9069 ( .A(\sub_x_53/A[30] ), .B(n4966), .Z(n4767) );
  HS65_LH_NOR2AX3 U9070 ( .A(n4535), .B(n5152), .Z(n6121) );
  HS65_LH_NAND2X2 U9071 ( .A(n4551), .B(n4550), .Z(n4580) );
  HS65_LH_NAND2X2 U9072 ( .A(n5217), .B(n4563), .Z(n4564) );
  HS65_LLS_XNOR2X3 U9073 ( .A(n4577), .B(n4576), .Z(n4605) );
  HS65_LH_CBI4I1X3 U9074 ( .A(n5648), .B(n5321), .C(n4804), .D(\lte_x_59/B[3] ), .Z(n4586) );
  HS65_LH_OAI222X2 U9075 ( .A(n4796), .B(n4583), .C(n2848), .D(n4582), .E(
        n2893), .F(n5041), .Z(n4584) );
  HS65_LHS_XNOR2X3 U9076 ( .A(\lte_x_59/B[3] ), .B(n5321), .Z(n4763) );
  HS65_LH_AOI22X1 U9077 ( .A(\lte_x_59/B[7] ), .B(n4588), .C(n4587), .D(
        \lte_x_59/B[8] ), .Z(n4589) );
  HS65_LH_CBI4I1X3 U9078 ( .A(n3582), .B(n5030), .C(n5647), .D(\lte_x_59/B[7] ), .Z(n4612) );
  HS65_LH_CNIVX3 U9079 ( .A(n4638), .Z(n4639) );
  HS65_LH_NAND2X5 U9080 ( .A(n5032), .B(n4796), .Z(n5322) );
  HS65_LH_CB4I1X9 U9081 ( .A(n4657), .B(n8495), .C(n4656), .D(n5041), .Z(n5388) );
  HS65_LH_NAND2X7 U9083 ( .A(n4711), .B(n4976), .Z(n5564) );
  HS65_LH_NAND2X7 U9084 ( .A(n4725), .B(n5422), .Z(n5286) );
  HS65_LH_NAND4ABX3 U9085 ( .A(n5426), .B(n5571), .C(n5286), .D(n5289), .Z(
        n4691) );
  HS65_LH_NAND3X2 U9086 ( .A(n3384), .B(n2853), .C(n5564), .Z(n4723) );
  HS65_LH_NOR3X1 U9087 ( .A(n4713), .B(n8833), .C(n4712), .Z(n4719) );
  HS65_LH_OAI31X1 U9088 ( .A(n4717), .B(n8427), .C(n7868), .D(n4716), .Z(n4718) );
  HS65_LHS_XNOR2X3 U9089 ( .A(\lte_x_59/B[9] ), .B(n5053), .Z(n4870) );
  HS65_LHS_XNOR2X3 U9090 ( .A(n5061), .B(\lte_x_59/B[14] ), .Z(n4945) );
  HS65_LHS_XNOR2X3 U9091 ( .A(\lte_x_59/B[24] ), .B(n5180), .Z(n5188) );
  HS65_LH_NOR3X4 U9092 ( .A(n4815), .B(n4814), .C(n4813), .Z(n4831) );
  HS65_LH_NAND3X2 U9093 ( .A(n5021), .B(n3582), .C(\lte_x_59/B[16] ), .Z(n4851) );
  HS65_LH_OAI21X3 U9094 ( .A(n4855), .B(n5204), .C(n4854), .Z(n4859) );
  HS65_LH_OAI21X3 U9095 ( .A(n4857), .B(n5656), .C(n4856), .Z(n4858) );
  HS65_LLS_XOR2X6 U9096 ( .A(n4864), .B(n5633), .Z(n4865) );
  HS65_LH_NAND2X7 U9097 ( .A(n7631), .B(n4865), .Z(n4866) );
  HS65_LH_OAI21X3 U9098 ( .A(n4870), .B(n5656), .C(n4869), .Z(n4871) );
  HS65_LH_CBI4I1X3 U9099 ( .A(n5648), .B(n5053), .C(n5647), .D(\lte_x_59/B[9] ), .Z(n4890) );
  HS65_LH_CBI4I1X3 U9100 ( .A(n5648), .B(n5061), .C(n3443), .D(
        \lte_x_59/B[14] ), .Z(n4940) );
  HS65_LH_NAND2X2 U9101 ( .A(\lte_x_59/B[24] ), .B(n3382), .Z(n5442) );
  HS65_LH_CBI4I1X3 U9102 ( .A(n5009), .B(n5586), .C(n5585), .D(n5115), .Z(
        n4978) );
  HS65_LH_NOR3AX2 U9103 ( .A(n5022), .B(n5023), .C(n4985), .Z(n4987) );
  HS65_LH_NOR2X3 U9104 ( .A(n5041), .B(n5040), .Z(n5042) );
  HS65_LH_NOR2X2 U9105 ( .A(n4796), .B(n5032), .Z(n5033) );
  HS65_LH_NOR2X2 U9106 ( .A(n5088), .B(n5130), .Z(n5036) );
  HS65_LH_OAI21X3 U9107 ( .A(n5322), .B(n5042), .C(n5328), .Z(n5098) );
  HS65_LH_AND2X4 U9109 ( .A(n5126), .B(n5125), .Z(n5155) );
  HS65_LH_CBI4I1X3 U9110 ( .A(n5648), .B(n5136), .C(n3443), .D(\sub_x_53/A[0] ), .Z(n5137) );
  HS65_LH_NAND2X7 U9111 ( .A(n5168), .B(n5167), .Z(n5695) );
  HS65_LHS_XOR2X3 U9112 ( .A(n5696), .B(n5695), .Z(n5169) );
  HS65_LH_CBI4I1X3 U9113 ( .A(n5648), .B(n5180), .C(n5647), .D(
        \lte_x_59/B[24] ), .Z(n5181) );
  HS65_LH_NAND3X3 U9116 ( .A(n5292), .B(n5362), .C(n5291), .Z(n5354) );
  HS65_LH_NOR2X2 U9118 ( .A(n5321), .B(n5320), .Z(n5323) );
  HS65_LH_AOI21X2 U9119 ( .A(n5433), .B(n5432), .C(n5431), .Z(n5440) );
  HS65_LH_NAND2X2 U9120 ( .A(\lte_x_59/B[21] ), .B(n3377), .Z(n5434) );
  HS65_LH_NAND2X2 U9121 ( .A(\lte_x_59/B[22] ), .B(n2869), .Z(n5435) );
  HS65_LH_AOI21X2 U9122 ( .A(n5438), .B(n5437), .C(n5436), .Z(n5439) );
  HS65_LL_AOI12X2 U9123 ( .A(n5495), .B(n5494), .C(n5493), .Z(n5496) );
  HS65_LH_NAND3X5 U9124 ( .A(n5574), .B(n5582), .C(n5562), .Z(n5527) );
  HS65_LH_NAND4ABX3 U9125 ( .A(n5512), .B(n5511), .C(n5529), .D(n5536), .Z(
        n5513) );
  HS65_LL_NAND4ABX3 U9126 ( .A(n5558), .B(n5557), .C(n5556), .D(n5555), .Z(
        n5560) );
  HS65_LH_OAI21X3 U9127 ( .A(n5578), .B(n5577), .C(n5576), .Z(n5579) );
  HS65_LHS_XNOR2X3 U9128 ( .A(\lte_x_59/B[22] ), .B(n5654), .Z(n5655) );
  HS65_LHS_XNOR2X3 U9129 ( .A(n5697), .B(n7118), .Z(n5698) );
  HS65_LL_AOI22X1 U9130 ( .A(n8868), .B(n9032), .C(n9369), .D(n9047), .Z(n7858) );
  HS65_LH_AND2X4 U9131 ( .A(n5850), .B(n5717), .Z(\u_DataPath/toPC2_i [0]) );
  HS65_LH_CNIVX3 U9132 ( .A(n5748), .Z(n5749) );
  HS65_LH_CNIVX3 U9133 ( .A(n5767), .Z(n5768) );
  HS65_LH_CNIVX3 U9134 ( .A(n5817), .Z(n5818) );
  HS65_LH_AOI21X2 U9136 ( .A(n5890), .B(n5892), .C(n6042), .Z(n5841) );
  HS65_LHS_XOR2X3 U9137 ( .A(n5850), .B(n5849), .Z(\u_DataPath/toPC2_i [1]) );
  HS65_LH_OR2X4 U9138 ( .A(n9341), .B(n9202), .Z(n5851) );
  HS65_LLS_XNOR2X3 U9139 ( .A(n5857), .B(n5856), .Z(\u_DataPath/toPC2_i [31])
         );
  HS65_LHS_XNOR2X3 U9140 ( .A(n5905), .B(n5904), .Z(\u_DataPath/toPC2_i [21])
         );
  HS65_LH_AND2X4 U9141 ( .A(n6049), .B(n5918), .Z(
        \u_DataPath/u_execute/resAdd1_i [0]) );
  HS65_LH_CNIVX3 U9145 ( .A(n5971), .Z(n5972) );
  HS65_LH_CNIVX3 U9146 ( .A(n5995), .Z(n5996) );
  HS65_LH_CNIVX3 U9147 ( .A(n5998), .Z(n6002) );
  HS65_LH_CNIVX3 U9148 ( .A(n6026), .Z(n6027) );
  HS65_LH_AOI21X2 U9149 ( .A(n5890), .B(n6095), .C(n6042), .Z(n6043) );
  HS65_LHS_XOR2X3 U9150 ( .A(n6049), .B(n6048), .Z(
        \u_DataPath/u_execute/resAdd1_i [1]) );
  HS65_LH_NAND2X2 U9152 ( .A(n6099), .B(n6098), .Z(n6104) );
  HS65_LHS_XNOR2X3 U9153 ( .A(n6108), .B(n6107), .Z(
        \u_DataPath/u_execute/resAdd1_i [24]) );
  HS65_LHS_XNOR2X3 U9154 ( .A(n6112), .B(n6111), .Z(
        \u_DataPath/u_execute/resAdd1_i [22]) );
  HS65_LH_AOI22X1 U9155 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][30] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][30] ), .D(
        n6362), .Z(n6130) );
  HS65_LH_BFX9 U9156 ( .A(n6162), .Z(n7265) );
  HS65_LH_NOR2X6 U9157 ( .A(n6150), .B(n6151), .Z(n6363) );
  HS65_LH_NOR4ABX2 U9158 ( .A(n6130), .B(n6129), .C(n6128), .D(n6127), .Z(
        n6161) );
  HS65_LH_BFX9 U9159 ( .A(n6370), .Z(n7165) );
  HS65_LH_BFX9 U9160 ( .A(n6371), .Z(n7273) );
  HS65_LH_NOR2X13 U9161 ( .A(n6150), .B(n6133), .Z(n6628) );
  HS65_LH_NOR4ABX2 U9162 ( .A(n6137), .B(n6136), .C(n6135), .D(n6134), .Z(
        n6160) );
  HS65_LH_NOR2X6 U9163 ( .A(n6148), .B(n6139), .Z(n6377) );
  HS65_LH_NAND4ABX3 U9164 ( .A(n6144), .B(n6143), .C(n6142), .D(n6141), .Z(
        n6159) );
  HS65_LH_BFX9 U9165 ( .A(n6383), .Z(n7292) );
  HS65_LH_NOR2X6 U9166 ( .A(n6150), .B(n6152), .Z(n7295) );
  HS65_LH_NOR2X6 U9167 ( .A(n6153), .B(n6151), .Z(n6385) );
  HS65_LH_NAND4ABX3 U9168 ( .A(n6157), .B(n6156), .C(n6155), .D(n6154), .Z(
        n6158) );
  HS65_LH_AOI22X1 U9169 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][16] ), .D(
        n6362), .Z(n6166) );
  HS65_LH_AO22X9 U9170 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][16] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][16] ), .D(
        n9371), .Z(n6164) );
  HS65_LH_NOR4ABX2 U9171 ( .A(n6166), .B(n6165), .C(n6164), .D(n6163), .Z(
        n6184) );
  HS65_LH_NOR4ABX2 U9172 ( .A(n6170), .B(n6169), .C(n6168), .D(n6167), .Z(
        n6183) );
  HS65_LH_NAND4ABX3 U9173 ( .A(n6176), .B(n6175), .C(n6174), .D(n6173), .Z(
        n6182) );
  HS65_LH_AO22X9 U9174 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][16] ), .B(n6317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][16] ), .D(
        n7292), .Z(n6179) );
  HS65_LH_AOI22X1 U9175 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][16] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ), .D(
        n6384), .Z(n6178) );
  HS65_LH_NAND4ABX3 U9176 ( .A(n6180), .B(n6179), .C(n6178), .D(n6177), .Z(
        n6181) );
  HS65_LH_NOR4ABX2 U9177 ( .A(n6188), .B(n6187), .C(n6186), .D(n6185), .Z(
        n6204) );
  HS65_LH_NOR4ABX2 U9178 ( .A(n6192), .B(n6191), .C(n6190), .D(n6189), .Z(
        n6203) );
  HS65_LH_NAND4ABX3 U9179 ( .A(n6196), .B(n6195), .C(n6194), .D(n6193), .Z(
        n6202) );
  HS65_LH_AOI22X1 U9180 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][21] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ), .D(
        n6384), .Z(n6198) );
  HS65_LH_NAND4ABX3 U9181 ( .A(n6200), .B(n6199), .C(n6198), .D(n6197), .Z(
        n6201) );
  HS65_LH_AO22X9 U9182 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][27] ), .D(
        n9371), .Z(n6206) );
  HS65_LH_NOR4ABX2 U9183 ( .A(n6208), .B(n6207), .C(n6206), .D(n6205), .Z(
        n6224) );
  HS65_LH_NOR4ABX2 U9184 ( .A(n6212), .B(n6211), .C(n6210), .D(n6209), .Z(
        n6223) );
  HS65_LH_NAND4ABX3 U9185 ( .A(n6216), .B(n6215), .C(n6214), .D(n6213), .Z(
        n6222) );
  HS65_LH_AOI22X1 U9186 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][27] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][27] ), .D(
        n6384), .Z(n6218) );
  HS65_LH_NAND4ABX3 U9187 ( .A(n6220), .B(n6219), .C(n6218), .D(n6217), .Z(
        n6221) );
  HS65_LH_AO22X9 U9188 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][23] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][23] ), .D(
        n9372), .Z(n6226) );
  HS65_LH_NOR4ABX2 U9189 ( .A(n6228), .B(n6227), .C(n6226), .D(n6225), .Z(
        n6244) );
  HS65_LH_NOR4ABX2 U9190 ( .A(n6232), .B(n6231), .C(n6230), .D(n6229), .Z(
        n6243) );
  HS65_LH_NAND4ABX3 U9191 ( .A(n6236), .B(n6235), .C(n6234), .D(n6233), .Z(
        n6242) );
  HS65_LH_BFX9 U9192 ( .A(n6317), .Z(n7293) );
  HS65_LH_AOI22X1 U9193 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][23] ), .D(
        n6384), .Z(n6238) );
  HS65_LH_NAND4ABX3 U9194 ( .A(n6240), .B(n6239), .C(n6238), .D(n6237), .Z(
        n6241) );
  HS65_LH_AO22X9 U9195 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][11] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][11] ), .D(
        n9372), .Z(n6246) );
  HS65_LH_NOR4ABX2 U9196 ( .A(n6248), .B(n6247), .C(n6246), .D(n6245), .Z(
        n6264) );
  HS65_LH_NOR4ABX2 U9197 ( .A(n6252), .B(n6251), .C(n6250), .D(n6249), .Z(
        n6263) );
  HS65_LH_NAND4ABX3 U9198 ( .A(n6256), .B(n6255), .C(n6254), .D(n6253), .Z(
        n6262) );
  HS65_LH_AOI22X1 U9199 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][11] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][11] ), .D(
        n6384), .Z(n6258) );
  HS65_LH_NAND4ABX3 U9200 ( .A(n6260), .B(n6259), .C(n6258), .D(n6257), .Z(
        n6261) );
  HS65_LH_AOI22X1 U9201 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][22] ), .B(n6617), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][22] ), .D(
        n6362), .Z(n6268) );
  HS65_LH_NOR4ABX2 U9202 ( .A(n6268), .B(n6267), .C(n6266), .D(n6265), .Z(
        n6284) );
  HS65_LH_NOR4ABX2 U9203 ( .A(n6272), .B(n6271), .C(n6270), .D(n6269), .Z(
        n6283) );
  HS65_LH_NAND4ABX3 U9204 ( .A(n6276), .B(n6275), .C(n6274), .D(n6273), .Z(
        n6282) );
  HS65_LH_AOI22X1 U9205 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][22] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][22] ), .D(
        n6384), .Z(n6278) );
  HS65_LH_NAND4ABX3 U9206 ( .A(n6280), .B(n6279), .C(n6278), .D(n6277), .Z(
        n6281) );
  HS65_LH_NOR4ABX2 U9207 ( .A(n6288), .B(n6287), .C(n6286), .D(n6285), .Z(
        n6304) );
  HS65_LH_NOR4ABX2 U9208 ( .A(n6292), .B(n6291), .C(n6290), .D(n6289), .Z(
        n6303) );
  HS65_LH_NAND4ABX3 U9209 ( .A(n6296), .B(n6295), .C(n6294), .D(n6293), .Z(
        n6302) );
  HS65_LH_AOI22X1 U9210 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][24] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ), .D(
        n6384), .Z(n6298) );
  HS65_LH_NAND4ABX3 U9211 ( .A(n6300), .B(n6299), .C(n6298), .D(n6297), .Z(
        n6301) );
  HS65_LH_NOR4ABX2 U9212 ( .A(n6308), .B(n6307), .C(n6306), .D(n6305), .Z(
        n6325) );
  HS65_LH_NOR4ABX2 U9213 ( .A(n6312), .B(n6311), .C(n6310), .D(n6309), .Z(
        n6324) );
  HS65_LH_NAND4ABX3 U9214 ( .A(n6316), .B(n6315), .C(n6314), .D(n6313), .Z(
        n6323) );
  HS65_LH_AOI22X1 U9215 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][14] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][14] ), .D(
        n6384), .Z(n6319) );
  HS65_LH_NAND4ABX3 U9216 ( .A(n6321), .B(n6320), .C(n6319), .D(n6318), .Z(
        n6322) );
  HS65_LH_NAND3X5 U9217 ( .A(\u_DataPath/jaddr_i [19]), .B(
        \u_DataPath/jaddr_i [18]), .C(n2881), .Z(n6334) );
  HS65_LH_NOR2X6 U9218 ( .A(\u_DataPath/jaddr_i [19]), .B(n8184), .Z(n6340) );
  HS65_LH_NOR4ABX2 U9220 ( .A(n6330), .B(n6329), .C(n6328), .D(n6327), .Z(
        n6361) );
  HS65_LH_NOR2X6 U9221 ( .A(n6353), .B(n6332), .Z(n6957) );
  HS65_LH_AOI22X1 U9222 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][18] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][18] ), .D(
        n6957), .Z(n6337) );
  HS65_LH_BFX9 U9223 ( .A(n6747), .Z(n7517) );
  HS65_LH_NOR2X6 U9224 ( .A(n6350), .B(n6333), .Z(n6675) );
  HS65_LH_NOR2X6 U9225 ( .A(n6350), .B(n6334), .Z(n7319) );
  HS65_LH_NOR4ABX2 U9226 ( .A(n6338), .B(n6337), .C(n6336), .D(n6335), .Z(
        n6360) );
  HS65_LH_NAND2X7 U9227 ( .A(\u_DataPath/jaddr_i [20]), .B(n6340), .Z(n6342)
         );
  HS65_LH_AO22X9 U9228 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][18] ), .B(n7522), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][18] ), .Z(n6346)
         );
  HS65_LH_NOR2X6 U9230 ( .A(n6353), .B(n6342), .Z(n6753) );
  HS65_LH_NOR2X6 U9231 ( .A(n6349), .B(n6342), .Z(n6684) );
  HS65_LH_NAND4ABX3 U9232 ( .A(n6346), .B(n6345), .C(n6344), .D(n6343), .Z(
        n6359) );
  HS65_LH_NAND2X7 U9233 ( .A(n8184), .B(n6347), .Z(n6351) );
  HS65_LH_NOR2X6 U9234 ( .A(n6348), .B(n6351), .Z(n7330) );
  HS65_LH_NOR2X6 U9235 ( .A(n6349), .B(n6351), .Z(n7329) );
  HS65_LH_NAND2X7 U9236 ( .A(\u_DataPath/jaddr_i [18]), .B(n6347), .Z(n6352)
         );
  HS65_LH_NOR2X6 U9237 ( .A(n6348), .B(n6352), .Z(n7332) );
  HS65_LH_NOR2X6 U9238 ( .A(n6350), .B(n6351), .Z(n7331) );
  HS65_LH_NOR2X6 U9239 ( .A(n6353), .B(n6351), .Z(n6690) );
  HS65_LH_NAND4ABX3 U9240 ( .A(n6357), .B(n6356), .C(n6355), .D(n6354), .Z(
        n6358) );
  HS65_LH_BFX9 U9241 ( .A(n6617), .Z(n6595) );
  HS65_LH_BFX9 U9242 ( .A(n6362), .Z(n7264) );
  HS65_LH_AO22X9 U9243 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][15] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][15] ), .D(
        n7266), .Z(n6367) );
  HS65_LH_AO22X9 U9244 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][15] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][15] ), .D(
        n7267), .Z(n6366) );
  HS65_LH_NOR4ABX2 U9245 ( .A(n6369), .B(n6368), .C(n6367), .D(n6366), .Z(
        n6393) );
  HS65_LH_AO22X9 U9247 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][15] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][15] ), .D(
        n7274), .Z(n6373) );
  HS65_LH_NOR4ABX2 U9248 ( .A(n6375), .B(n6374), .C(n6373), .D(n6372), .Z(
        n6392) );
  HS65_LH_NAND4ABX3 U9249 ( .A(n6381), .B(n6380), .C(n6379), .D(n6378), .Z(
        n6391) );
  HS65_LH_AO22X9 U9250 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][15] ), .D(
        n7291), .Z(n6389) );
  HS65_LH_BFX9 U9251 ( .A(n6384), .Z(n7294) );
  HS65_LH_NAND4ABX3 U9252 ( .A(n6389), .B(n6388), .C(n6387), .D(n6386), .Z(
        n6390) );
  HS65_LH_AO22X9 U9253 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][10] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][10] ), .D(
        n7266), .Z(n6395) );
  HS65_LH_AO22X9 U9254 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][10] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][10] ), .D(
        n7267), .Z(n6394) );
  HS65_LH_NOR4ABX2 U9255 ( .A(n6397), .B(n6396), .C(n6395), .D(n6394), .Z(
        n6413) );
  HS65_LH_AO22X9 U9256 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][10] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][10] ), .D(
        n7274), .Z(n6399) );
  HS65_LH_NOR4ABX2 U9257 ( .A(n6401), .B(n6400), .C(n6399), .D(n6398), .Z(
        n6412) );
  HS65_LH_NAND4ABX3 U9258 ( .A(n6405), .B(n6404), .C(n6403), .D(n6402), .Z(
        n6411) );
  HS65_LH_NAND4ABX3 U9260 ( .A(n6409), .B(n6408), .C(n6407), .D(n6406), .Z(
        n6410) );
  HS65_LH_AO22X9 U9261 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][0] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ), .D(n7266), .Z(n6415) );
  HS65_LH_AO22X9 U9262 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][0] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][0] ), .D(n7267), .Z(n6414) );
  HS65_LH_NOR4ABX2 U9263 ( .A(n6417), .B(n6416), .C(n6415), .D(n6414), .Z(
        n6434) );
  HS65_LH_AOI22X1 U9264 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][0] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ), .D(
        n6600), .Z(n6421) );
  HS65_LH_AO22X9 U9265 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][0] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][0] ), .D(
        n7274), .Z(n6419) );
  HS65_LH_NOR4ABX2 U9266 ( .A(n6421), .B(n6420), .C(n6419), .D(n6418), .Z(
        n6433) );
  HS65_LH_NAND4ABX3 U9267 ( .A(n6425), .B(n6424), .C(n6423), .D(n6422), .Z(
        n6432) );
  HS65_LH_AOI22X3 U9269 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][0] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][0] ), .D(n7294), .Z(n6428) );
  HS65_LH_NAND4ABX3 U9270 ( .A(n6430), .B(n6429), .C(n6428), .D(n6427), .Z(
        n6431) );
  HS65_LH_AO22X9 U9271 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][7] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][7] ), .D(n7266), .Z(n6436) );
  HS65_LH_NOR4ABX2 U9273 ( .A(n6438), .B(n6437), .C(n6436), .D(n6435), .Z(
        n6454) );
  HS65_LH_AO22X9 U9274 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][7] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][7] ), .D(
        n7274), .Z(n6440) );
  HS65_LH_NOR4ABX2 U9275 ( .A(n6442), .B(n6441), .C(n6440), .D(n6439), .Z(
        n6453) );
  HS65_LH_NAND4ABX3 U9276 ( .A(n6446), .B(n6445), .C(n6444), .D(n6443), .Z(
        n6452) );
  HS65_LH_AOI22X3 U9278 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][7] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][7] ), .D(n7294), .Z(n6448) );
  HS65_LH_NAND4ABX3 U9279 ( .A(n6450), .B(n6449), .C(n6448), .D(n6447), .Z(
        n6451) );
  HS65_LH_AO22X9 U9280 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][8] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][8] ), .D(n7266), .Z(n6456) );
  HS65_LH_NOR4ABX2 U9282 ( .A(n6458), .B(n6457), .C(n6456), .D(n6455), .Z(
        n6474) );
  HS65_LH_AOI22X1 U9283 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][8] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][8] ), .D(
        n6600), .Z(n6462) );
  HS65_LH_AO22X9 U9284 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][8] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][8] ), .D(
        n7274), .Z(n6460) );
  HS65_LH_NOR4ABX2 U9285 ( .A(n6462), .B(n6461), .C(n6460), .D(n6459), .Z(
        n6473) );
  HS65_LH_NAND4ABX3 U9286 ( .A(n6466), .B(n6465), .C(n6464), .D(n6463), .Z(
        n6472) );
  HS65_LH_AO22X9 U9287 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][8] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][8] ), .D(n7291), .Z(n6470) );
  HS65_LH_AOI22X3 U9288 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][8] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][8] ), .D(n7294), .Z(n6468) );
  HS65_LH_NAND4ABX3 U9289 ( .A(n6470), .B(n6469), .C(n6468), .D(n6467), .Z(
        n6471) );
  HS65_LH_NOR4ABX2 U9290 ( .A(n6478), .B(n6477), .C(n6476), .D(n6475), .Z(
        n6494) );
  HS65_LH_AOI22X1 U9291 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][6] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][6] ), .D(
        n6600), .Z(n6482) );
  HS65_LH_NOR4ABX2 U9292 ( .A(n6482), .B(n6481), .C(n6480), .D(n6479), .Z(
        n6493) );
  HS65_LH_NAND4ABX3 U9293 ( .A(n6486), .B(n6485), .C(n6484), .D(n6483), .Z(
        n6492) );
  HS65_LH_NAND4ABX3 U9294 ( .A(n6490), .B(n6489), .C(n6488), .D(n6487), .Z(
        n6491) );
  HS65_LH_AO22X9 U9295 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][26] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][26] ), .D(
        n7266), .Z(n6496) );
  HS65_LH_AO22X9 U9296 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][26] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][26] ), .D(
        n7267), .Z(n6495) );
  HS65_LH_NOR4ABX2 U9297 ( .A(n6498), .B(n6497), .C(n6496), .D(n6495), .Z(
        n6514) );
  HS65_LH_AO22X9 U9298 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][26] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][26] ), .D(
        n7274), .Z(n6500) );
  HS65_LH_NOR4ABX2 U9299 ( .A(n6502), .B(n6501), .C(n6500), .D(n6499), .Z(
        n6513) );
  HS65_LH_NAND4ABX3 U9300 ( .A(n6506), .B(n6505), .C(n6504), .D(n6503), .Z(
        n6512) );
  HS65_LH_AO22X9 U9301 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][26] ), .D(
        n7291), .Z(n6510) );
  HS65_LH_AOI22X3 U9302 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][26] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][26] ), .D(
        n7294), .Z(n6508) );
  HS65_LH_NAND4ABX3 U9303 ( .A(n6510), .B(n6509), .C(n6508), .D(n6507), .Z(
        n6511) );
  HS65_LH_AO22X9 U9304 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][19] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ), .D(
        n7266), .Z(n6516) );
  HS65_LH_NOR4ABX2 U9306 ( .A(n6518), .B(n6517), .C(n6516), .D(n6515), .Z(
        n6534) );
  HS65_LH_AO22X9 U9307 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][19] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][19] ), .D(
        n7274), .Z(n6520) );
  HS65_LH_NOR4ABX2 U9308 ( .A(n6522), .B(n6521), .C(n6520), .D(n6519), .Z(
        n6533) );
  HS65_LH_NAND4ABX3 U9309 ( .A(n6526), .B(n6525), .C(n6524), .D(n6523), .Z(
        n6532) );
  HS65_LH_AO22X9 U9310 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][19] ), .D(
        n7291), .Z(n6530) );
  HS65_LH_AOI22X3 U9311 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][19] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][19] ), .D(
        n7294), .Z(n6528) );
  HS65_LH_NAND4ABX3 U9312 ( .A(n6530), .B(n6529), .C(n6528), .D(n6527), .Z(
        n6531) );
  HS65_LH_AO22X9 U9313 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][12] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][12] ), .D(
        n7266), .Z(n6536) );
  HS65_LH_NOR4ABX2 U9315 ( .A(n6538), .B(n6537), .C(n6536), .D(n6535), .Z(
        n6554) );
  HS65_LH_AO22X9 U9316 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][12] ), .D(
        n7274), .Z(n6540) );
  HS65_LH_NOR4ABX2 U9317 ( .A(n6542), .B(n6541), .C(n6540), .D(n6539), .Z(
        n6553) );
  HS65_LH_NAND4ABX3 U9318 ( .A(n6546), .B(n6545), .C(n6544), .D(n6543), .Z(
        n6552) );
  HS65_LH_AOI22X3 U9320 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][12] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][12] ), .D(
        n7294), .Z(n6548) );
  HS65_LH_NAND4ABX3 U9321 ( .A(n6550), .B(n6549), .C(n6548), .D(n6547), .Z(
        n6551) );
  HS65_LH_AO22X9 U9322 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][2] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][2] ), .D(n9371), .Z(n6556) );
  HS65_LH_NOR4ABX2 U9324 ( .A(n6558), .B(n6557), .C(n6556), .D(n6555), .Z(
        n6574) );
  HS65_LH_AOI22X1 U9325 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][2] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][2] ), .D(
        n6600), .Z(n6562) );
  HS65_LH_AO22X9 U9326 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][2] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][2] ), .D(
        n6627), .Z(n6560) );
  HS65_LH_AO22X9 U9327 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][2] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][2] ), .D(
        n6629), .Z(n6559) );
  HS65_LH_NOR4ABX2 U9328 ( .A(n6562), .B(n6561), .C(n6560), .D(n6559), .Z(
        n6573) );
  HS65_LH_NAND4ABX3 U9329 ( .A(n6566), .B(n6565), .C(n6564), .D(n6563), .Z(
        n6572) );
  HS65_LH_AO22X9 U9330 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][2] ), .D(n7291), .Z(n6570) );
  HS65_LH_AOI22X3 U9331 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][2] ), .D(n7294), .Z(n6568) );
  HS65_LH_NAND4ABX3 U9332 ( .A(n6570), .B(n6569), .C(n6568), .D(n6567), .Z(
        n6571) );
  HS65_LH_AO22X9 U9333 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][3] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][3] ), .D(n7266), .Z(n6576) );
  HS65_LH_AO22X9 U9334 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][3] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ), .D(n7267), .Z(n6575) );
  HS65_LH_NOR4ABX2 U9335 ( .A(n6578), .B(n6577), .C(n6576), .D(n6575), .Z(
        n6594) );
  HS65_LH_NOR4ABX2 U9336 ( .A(n6582), .B(n6581), .C(n6580), .D(n6579), .Z(
        n6593) );
  HS65_LH_NAND4ABX3 U9337 ( .A(n6586), .B(n6585), .C(n6584), .D(n6583), .Z(
        n6592) );
  HS65_LH_AO22X9 U9338 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][3] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][3] ), .D(n7291), .Z(n6590) );
  HS65_LH_AOI22X3 U9339 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][3] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][3] ), .D(n7294), .Z(n6588) );
  HS65_LH_NAND4ABX3 U9340 ( .A(n6590), .B(n6589), .C(n6588), .D(n6587), .Z(
        n6591) );
  HS65_LH_AO22X9 U9341 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][1] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][1] ), .D(n6619), .Z(n6596) );
  HS65_LH_NOR4ABX2 U9342 ( .A(n6599), .B(n6598), .C(n6597), .D(n6596), .Z(
        n6616) );
  HS65_LH_AO22X9 U9343 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][1] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][1] ), .D(
        n6629), .Z(n6601) );
  HS65_LH_NOR4ABX2 U9344 ( .A(n6604), .B(n6603), .C(n6602), .D(n6601), .Z(
        n6615) );
  HS65_LH_NAND4ABX3 U9345 ( .A(n6608), .B(n6607), .C(n6606), .D(n6605), .Z(
        n6614) );
  HS65_LH_AO22X9 U9346 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][1] ), .D(n7291), .Z(n6612) );
  HS65_LH_AOI22X3 U9347 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][1] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][1] ), .D(n7294), .Z(n6610) );
  HS65_LH_NAND4ABX3 U9348 ( .A(n6612), .B(n6611), .C(n6610), .D(n6609), .Z(
        n6613) );
  HS65_LH_BFX9 U9349 ( .A(n9370), .Z(n7266) );
  HS65_LH_AO22X9 U9350 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][4] ), .D(n7266), .Z(n6621) );
  HS65_LH_BFX9 U9351 ( .A(n6619), .Z(n7267) );
  HS65_LH_NOR4ABX2 U9353 ( .A(n6623), .B(n6622), .C(n6621), .D(n6620), .Z(
        n6649) );
  HS65_LH_BFX9 U9354 ( .A(n6626), .Z(n7275) );
  HS65_LH_AO22X9 U9355 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][4] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][4] ), .D(
        n7274), .Z(n6631) );
  HS65_LH_BFX9 U9356 ( .A(n6628), .Z(n7277) );
  HS65_LH_BFX9 U9357 ( .A(n6629), .Z(n7276) );
  HS65_LH_AO22X9 U9358 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][4] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][4] ), .D(
        n7276), .Z(n6630) );
  HS65_LH_NOR4ABX2 U9359 ( .A(n6633), .B(n6632), .C(n6631), .D(n6630), .Z(
        n6648) );
  HS65_LH_NAND4ABX3 U9360 ( .A(n6641), .B(n6640), .C(n6639), .D(n6638), .Z(
        n6647) );
  HS65_LH_NAND4ABX3 U9362 ( .A(n6645), .B(n6644), .C(n6643), .D(n6642), .Z(
        n6646) );
  HS65_LH_AO22X9 U9363 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][18] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][18] ), .D(
        n7266), .Z(n6651) );
  HS65_LH_AO22X9 U9364 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][18] ), .D(
        n7267), .Z(n6650) );
  HS65_LH_NOR4ABX2 U9365 ( .A(n6653), .B(n6652), .C(n6651), .D(n6650), .Z(
        n6669) );
  HS65_LH_AO22X9 U9367 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][18] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][18] ), .D(
        n7276), .Z(n6654) );
  HS65_LH_NOR4ABX2 U9368 ( .A(n6657), .B(n6656), .C(n6655), .D(n6654), .Z(
        n6668) );
  HS65_LH_NAND4ABX3 U9369 ( .A(n6661), .B(n6660), .C(n6659), .D(n6658), .Z(
        n6667) );
  HS65_LH_AOI22X3 U9370 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][18] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][18] ), .D(
        n7294), .Z(n6663) );
  HS65_LH_NAND4ABX3 U9371 ( .A(n6665), .B(n6664), .C(n6663), .D(n6662), .Z(
        n6666) );
  HS65_LH_NOR4ABX2 U9372 ( .A(n6674), .B(n6673), .C(n6672), .D(n6671), .Z(
        n6698) );
  HS65_LH_NOR4ABX2 U9373 ( .A(n6679), .B(n6678), .C(n6677), .D(n6676), .Z(
        n6697) );
  HS65_LH_BFX9 U9374 ( .A(n6752), .Z(n7439) );
  HS65_LH_NAND4ABX3 U9375 ( .A(n6688), .B(n6687), .C(n6686), .D(n6685), .Z(
        n6696) );
  HS65_LH_NAND4ABX3 U9376 ( .A(n6694), .B(n6693), .C(n6692), .D(n6691), .Z(
        n6695) );
  HS65_LH_NOR4ABX2 U9378 ( .A(n6702), .B(n6701), .C(n6700), .D(n6699), .Z(
        n6718) );
  HS65_LH_NOR4ABX2 U9379 ( .A(n6706), .B(n6705), .C(n6704), .D(n6703), .Z(
        n6717) );
  HS65_LH_NAND4ABX3 U9380 ( .A(n6710), .B(n6709), .C(n6708), .D(n6707), .Z(
        n6716) );
  HS65_LH_NAND4ABX3 U9381 ( .A(n6714), .B(n6713), .C(n6712), .D(n6711), .Z(
        n6715) );
  HS65_LH_NOR4ABX2 U9383 ( .A(n6722), .B(n6721), .C(n6720), .D(n6719), .Z(
        n6738) );
  HS65_LH_NOR4ABX2 U9384 ( .A(n6726), .B(n6725), .C(n6724), .D(n6723), .Z(
        n6737) );
  HS65_LH_NAND4ABX3 U9385 ( .A(n6730), .B(n6729), .C(n6728), .D(n6727), .Z(
        n6736) );
  HS65_LH_NAND4ABX3 U9386 ( .A(n6734), .B(n6733), .C(n6732), .D(n6731), .Z(
        n6735) );
  HS65_LH_NOR4ABX2 U9388 ( .A(n6744), .B(n6743), .C(n6742), .D(n6741), .Z(
        n6766) );
  HS65_LH_AOI22X1 U9389 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][19] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][19] ), .D(
        n6957), .Z(n6750) );
  HS65_LH_NOR4ABX2 U9390 ( .A(n6751), .B(n6750), .C(n6749), .D(n6748), .Z(
        n6765) );
  HS65_LH_NAND4ABX3 U9391 ( .A(n6758), .B(n6757), .C(n6756), .D(n6755), .Z(
        n6764) );
  HS65_LH_NAND4ABX3 U9392 ( .A(n6762), .B(n6761), .C(n6760), .D(n6759), .Z(
        n6763) );
  HS65_LH_NOR4ABX2 U9393 ( .A(n6770), .B(n6769), .C(n6768), .D(n6767), .Z(
        n6786) );
  HS65_LH_NOR4ABX2 U9394 ( .A(n6774), .B(n6773), .C(n6772), .D(n6771), .Z(
        n6785) );
  HS65_LH_NAND4ABX3 U9395 ( .A(n6778), .B(n6777), .C(n6776), .D(n6775), .Z(
        n6784) );
  HS65_LH_NAND4ABX3 U9396 ( .A(n6782), .B(n6781), .C(n6780), .D(n6779), .Z(
        n6783) );
  HS65_LL_NOR4ABX2 U9397 ( .A(n6786), .B(n6785), .C(n6784), .D(n6783), .Z(
        n8261) );
  HS65_LH_NOR4ABX2 U9398 ( .A(n6790), .B(n6789), .C(n6788), .D(n6787), .Z(
        n6806) );
  HS65_LH_NOR4ABX2 U9399 ( .A(n6794), .B(n6793), .C(n6792), .D(n6791), .Z(
        n6805) );
  HS65_LH_NAND4ABX3 U9400 ( .A(n6798), .B(n6797), .C(n6796), .D(n6795), .Z(
        n6804) );
  HS65_LH_NAND4ABX3 U9401 ( .A(n6802), .B(n6801), .C(n6800), .D(n6799), .Z(
        n6803) );
  HS65_LH_NOR4ABX2 U9402 ( .A(n6810), .B(n6809), .C(n6808), .D(n6807), .Z(
        n6826) );
  HS65_LH_NOR4ABX2 U9403 ( .A(n6814), .B(n6813), .C(n6812), .D(n6811), .Z(
        n6825) );
  HS65_LH_NAND4ABX3 U9404 ( .A(n6818), .B(n6817), .C(n6816), .D(n6815), .Z(
        n6824) );
  HS65_LH_NAND4ABX3 U9405 ( .A(n6822), .B(n6821), .C(n6820), .D(n6819), .Z(
        n6823) );
  HS65_LH_NOR4ABX2 U9407 ( .A(n6830), .B(n6829), .C(n6828), .D(n6827), .Z(
        n6846) );
  HS65_LH_NOR4ABX2 U9408 ( .A(n6834), .B(n6833), .C(n6832), .D(n6831), .Z(
        n6845) );
  HS65_LH_NAND4ABX3 U9409 ( .A(n6838), .B(n6837), .C(n6836), .D(n6835), .Z(
        n6844) );
  HS65_LH_NAND4ABX3 U9410 ( .A(n6842), .B(n6841), .C(n6840), .D(n6839), .Z(
        n6843) );
  HS65_LH_AO22X9 U9412 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][20] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][20] ), .D(
        n7267), .Z(n6847) );
  HS65_LH_NOR4ABX2 U9413 ( .A(n6850), .B(n6849), .C(n6848), .D(n6847), .Z(
        n6866) );
  HS65_LH_AO22X9 U9414 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][20] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][20] ), .D(
        n7274), .Z(n6852) );
  HS65_LH_NOR4ABX2 U9416 ( .A(n6854), .B(n6853), .C(n6852), .D(n6851), .Z(
        n6865) );
  HS65_LH_NAND4ABX3 U9417 ( .A(n6858), .B(n6857), .C(n6856), .D(n6855), .Z(
        n6864) );
  HS65_LH_AO22X9 U9418 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][20] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][20] ), .D(
        n7291), .Z(n6862) );
  HS65_LH_AOI22X3 U9419 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][20] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][20] ), .D(
        n7294), .Z(n6860) );
  HS65_LH_NAND4ABX3 U9420 ( .A(n6862), .B(n6861), .C(n6860), .D(n6859), .Z(
        n6863) );
  HS65_LH_AO22X9 U9421 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][31] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][31] ), .D(
        n7266), .Z(n6868) );
  HS65_LH_AO22X9 U9422 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][31] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][31] ), .D(
        n7267), .Z(n6867) );
  HS65_LH_NOR4ABX2 U9423 ( .A(n6870), .B(n6869), .C(n6868), .D(n6867), .Z(
        n6886) );
  HS65_LH_AOI22X1 U9424 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][31] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][31] ), .D(
        n6600), .Z(n6874) );
  HS65_LH_AO22X9 U9425 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][31] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][31] ), .D(
        n7274), .Z(n6872) );
  HS65_LH_AO22X9 U9426 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][31] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][31] ), .D(
        n7276), .Z(n6871) );
  HS65_LH_NOR4ABX2 U9427 ( .A(n6874), .B(n6873), .C(n6872), .D(n6871), .Z(
        n6885) );
  HS65_LH_NAND4ABX3 U9428 ( .A(n6878), .B(n6877), .C(n6876), .D(n6875), .Z(
        n6884) );
  HS65_LH_NAND4ABX3 U9429 ( .A(n6882), .B(n6881), .C(n6880), .D(n6879), .Z(
        n6883) );
  HS65_LH_AO22X9 U9430 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][17] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][17] ), .D(
        n7266), .Z(n6888) );
  HS65_LH_NOR4ABX2 U9432 ( .A(n6890), .B(n6889), .C(n6888), .D(n6887), .Z(
        n6906) );
  HS65_LH_AOI22X1 U9433 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][17] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][17] ), .D(
        n6600), .Z(n6894) );
  HS65_LH_AO22X9 U9434 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][17] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ), .D(
        n7274), .Z(n6892) );
  HS65_LH_AO22X9 U9435 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][17] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][17] ), .D(
        n7276), .Z(n6891) );
  HS65_LH_NOR4ABX2 U9436 ( .A(n6894), .B(n6893), .C(n6892), .D(n6891), .Z(
        n6905) );
  HS65_LH_NAND4ABX3 U9437 ( .A(n6898), .B(n6897), .C(n6896), .D(n6895), .Z(
        n6904) );
  HS65_LH_NAND4ABX3 U9439 ( .A(n6902), .B(n6901), .C(n6900), .D(n6899), .Z(
        n6903) );
  HS65_LH_AO22X9 U9440 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][28] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][28] ), .D(
        n7266), .Z(n6908) );
  HS65_LH_NOR4ABX2 U9442 ( .A(n6910), .B(n6909), .C(n6908), .D(n6907), .Z(
        n6926) );
  HS65_LH_AO22X9 U9443 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][28] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ), .D(
        n7274), .Z(n6912) );
  HS65_LH_AO22X9 U9444 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][28] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][28] ), .D(
        n7276), .Z(n6911) );
  HS65_LH_NOR4ABX2 U9445 ( .A(n6914), .B(n6913), .C(n6912), .D(n6911), .Z(
        n6925) );
  HS65_LH_NAND4ABX3 U9446 ( .A(n6918), .B(n6917), .C(n6916), .D(n6915), .Z(
        n6924) );
  HS65_LH_AO22X9 U9447 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][28] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][28] ), .D(
        n7291), .Z(n6922) );
  HS65_LH_AOI22X3 U9448 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][28] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][28] ), .D(
        n7294), .Z(n6920) );
  HS65_LH_NAND4ABX3 U9449 ( .A(n6922), .B(n6921), .C(n6920), .D(n6919), .Z(
        n6923) );
  HS65_LH_AO22X9 U9450 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][5] ), .D(n7266), .Z(n6930) );
  HS65_LH_AO22X9 U9451 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][5] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][5] ), .D(n7267), .Z(n6929) );
  HS65_LH_NOR4ABX2 U9452 ( .A(n6932), .B(n6931), .C(n6930), .D(n6929), .Z(
        n6950) );
  HS65_LH_AO22X9 U9453 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][5] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][5] ), .D(
        n7274), .Z(n6934) );
  HS65_LH_AO22X9 U9454 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][5] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][5] ), .D(
        n7276), .Z(n6933) );
  HS65_LH_NOR4ABX2 U9455 ( .A(n6936), .B(n6935), .C(n6934), .D(n6933), .Z(
        n6949) );
  HS65_LH_NAND4ABX3 U9456 ( .A(n6940), .B(n6939), .C(n6938), .D(n6937), .Z(
        n6948) );
  HS65_LH_AOI22X3 U9457 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][5] ), .D(n7294), .Z(n6944) );
  HS65_LH_NAND4ABX3 U9458 ( .A(n6946), .B(n6945), .C(n6944), .D(n6943), .Z(
        n6947) );
  HS65_LH_NOR4ABX2 U9459 ( .A(n6956), .B(n6955), .C(n6954), .D(n6953), .Z(
        n6975) );
  HS65_LH_NOR4ABX2 U9460 ( .A(n6961), .B(n6960), .C(n6959), .D(n6958), .Z(
        n6974) );
  HS65_LH_NAND4ABX3 U9461 ( .A(n6965), .B(n6964), .C(n6963), .D(n6962), .Z(
        n6973) );
  HS65_LH_NAND4ABX3 U9462 ( .A(n6971), .B(n6970), .C(n6969), .D(n6968), .Z(
        n6972) );
  HS65_LH_NOR4ABX2 U9463 ( .A(n6979), .B(n6978), .C(n6977), .D(n6976), .Z(
        n6995) );
  HS65_LH_AOI22X1 U9464 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][13] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][13] ), .D(
        n6957), .Z(n6982) );
  HS65_LH_NOR4ABX2 U9465 ( .A(n6983), .B(n6982), .C(n6981), .D(n6980), .Z(
        n6994) );
  HS65_LH_NAND4ABX3 U9466 ( .A(n6987), .B(n6986), .C(n6985), .D(n6984), .Z(
        n6993) );
  HS65_LH_NAND4ABX3 U9467 ( .A(n6991), .B(n6990), .C(n6989), .D(n6988), .Z(
        n6992) );
  HS65_LH_NOR4ABX2 U9468 ( .A(n6999), .B(n6998), .C(n6997), .D(n6996), .Z(
        n7015) );
  HS65_LH_AOI22X1 U9469 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][22] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][22] ), .D(
        n6957), .Z(n7002) );
  HS65_LH_NOR4ABX2 U9470 ( .A(n7003), .B(n7002), .C(n7001), .D(n7000), .Z(
        n7014) );
  HS65_LH_NAND4ABX3 U9471 ( .A(n7007), .B(n7006), .C(n7005), .D(n7004), .Z(
        n7013) );
  HS65_LH_NAND4ABX3 U9472 ( .A(n7011), .B(n7010), .C(n7009), .D(n7008), .Z(
        n7012) );
  HS65_LH_NOR4ABX2 U9473 ( .A(n7019), .B(n7018), .C(n7017), .D(n7016), .Z(
        n7035) );
  HS65_LH_AOI22X1 U9474 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][9] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ), .D(n6957), .Z(n7022) );
  HS65_LH_NOR4ABX2 U9475 ( .A(n7023), .B(n7022), .C(n7021), .D(n7020), .Z(
        n7034) );
  HS65_LH_NAND4ABX3 U9476 ( .A(n7027), .B(n7026), .C(n7025), .D(n7024), .Z(
        n7033) );
  HS65_LH_NAND4ABX3 U9477 ( .A(n7031), .B(n7030), .C(n7029), .D(n7028), .Z(
        n7032) );
  HS65_LH_NOR4ABX2 U9478 ( .A(n7039), .B(n7038), .C(n7037), .D(n7036), .Z(
        n7055) );
  HS65_LH_AOI22X1 U9479 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][25] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ), .D(
        n6957), .Z(n7042) );
  HS65_LH_NOR4ABX2 U9480 ( .A(n7043), .B(n7042), .C(n7041), .D(n7040), .Z(
        n7054) );
  HS65_LH_NAND4ABX3 U9481 ( .A(n7047), .B(n7046), .C(n7045), .D(n7044), .Z(
        n7053) );
  HS65_LH_NAND4ABX3 U9482 ( .A(n7051), .B(n7050), .C(n7049), .D(n7048), .Z(
        n7052) );
  HS65_LH_NOR4ABX2 U9483 ( .A(n7059), .B(n7058), .C(n7057), .D(n7056), .Z(
        n7075) );
  HS65_LH_AOI22X1 U9484 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][11] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][11] ), .D(
        n6957), .Z(n7062) );
  HS65_LH_NOR4ABX2 U9485 ( .A(n7063), .B(n7062), .C(n7061), .D(n7060), .Z(
        n7074) );
  HS65_LH_NAND4ABX3 U9486 ( .A(n7067), .B(n7066), .C(n7065), .D(n7064), .Z(
        n7073) );
  HS65_LH_NAND4ABX3 U9487 ( .A(n7071), .B(n7070), .C(n7069), .D(n7068), .Z(
        n7072) );
  HS65_LH_NOR2X6 U9488 ( .A(n7078), .B(n7077), .Z(n7082) );
  HS65_LH_NOR2X6 U9489 ( .A(n7080), .B(n7079), .Z(n7081) );
  HS65_LH_NAND2X7 U9491 ( .A(n7088), .B(n7087), .Z(n7093) );
  HS65_LH_NOR2X6 U9492 ( .A(\u_DataPath/cw_exmem_i [5]), .B(
        \u_DataPath/cw_exmem_i [3]), .Z(n7097) );
  HS65_LH_NAND2X7 U9493 ( .A(n7098), .B(n7097), .Z(n7114) );
  HS65_LH_NOR2X2 U9494 ( .A(n8426), .B(n9401), .Z(n8564) );
  HS65_LH_AO22X9 U9495 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][9] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][9] ), .D(n9371), .Z(n7124) );
  HS65_LH_NOR4ABX2 U9496 ( .A(n7126), .B(n7125), .C(n7124), .D(n7123), .Z(
        n7142) );
  HS65_LH_NOR4ABX2 U9498 ( .A(n7130), .B(n7129), .C(n7128), .D(n7127), .Z(
        n7141) );
  HS65_LH_NAND4ABX3 U9499 ( .A(n7134), .B(n7133), .C(n7132), .D(n7131), .Z(
        n7140) );
  HS65_LH_AOI22X1 U9501 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][9] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][9] ), .D(n7294), .Z(n7136) );
  HS65_LH_NAND4ABX3 U9502 ( .A(n7138), .B(n7137), .C(n7136), .D(n7135), .Z(
        n7139) );
  HS65_LH_NOR4ABX2 U9503 ( .A(n7142), .B(n7141), .C(n7140), .D(n7139), .Z(
        n8336) );
  HS65_LH_AO22X9 U9504 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][25] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][25] ), .D(
        n9372), .Z(n7144) );
  HS65_LH_NOR4ABX2 U9505 ( .A(n7146), .B(n7145), .C(n7144), .D(n7143), .Z(
        n7160) );
  HS65_LH_NOR4ABX2 U9507 ( .A(n7150), .B(n7149), .C(n7148), .D(n7147), .Z(
        n7159) );
  HS65_LH_AO22X9 U9508 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][25] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][25] ), .D(
        n7291), .Z(n7156) );
  HS65_LH_AOI22X1 U9509 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][25] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][25] ), .D(
        n6384), .Z(n7154) );
  HS65_LH_NAND4ABX3 U9510 ( .A(n7156), .B(n7155), .C(n7154), .D(n7153), .Z(
        n7157) );
  HS65_LH_NOR4ABX2 U9511 ( .A(n7160), .B(n7159), .C(n7158), .D(n7157), .Z(
        n8329) );
  HS65_LH_NOR4ABX2 U9512 ( .A(n7164), .B(n7163), .C(n7162), .D(n7161), .Z(
        n7183) );
  HS65_LH_NOR4ABX2 U9513 ( .A(n7169), .B(n7168), .C(n7167), .D(n7166), .Z(
        n7182) );
  HS65_LH_NAND4ABX3 U9514 ( .A(n7175), .B(n7174), .C(n7173), .D(n7172), .Z(
        n7181) );
  HS65_LH_AOI22X1 U9515 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][13] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][13] ), .D(
        n6384), .Z(n7177) );
  HS65_LH_NAND4ABX3 U9516 ( .A(n7179), .B(n7178), .C(n7177), .D(n7176), .Z(
        n7180) );
  HS65_LH_NOR4ABX2 U9517 ( .A(n7183), .B(n7182), .C(n7181), .D(n7180), .Z(
        n8342) );
  HS65_LH_NOR4ABX2 U9518 ( .A(n7187), .B(n7186), .C(n7185), .D(n7184), .Z(
        n7203) );
  HS65_LH_AOI22X1 U9519 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][15] ), .D(
        n6957), .Z(n7190) );
  HS65_LH_NOR4ABX2 U9520 ( .A(n7191), .B(n7190), .C(n7189), .D(n7188), .Z(
        n7202) );
  HS65_LH_NAND4ABX3 U9521 ( .A(n7195), .B(n7194), .C(n7193), .D(n7192), .Z(
        n7201) );
  HS65_LH_NAND4ABX3 U9522 ( .A(n7199), .B(n7198), .C(n7197), .D(n7196), .Z(
        n7200) );
  HS65_LH_NOR4ABX2 U9523 ( .A(n7207), .B(n7206), .C(n7205), .D(n7204), .Z(
        n7223) );
  HS65_LH_AOI22X1 U9524 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][10] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ), .D(
        n6957), .Z(n7210) );
  HS65_LH_NOR4ABX2 U9525 ( .A(n7211), .B(n7210), .C(n7209), .D(n7208), .Z(
        n7222) );
  HS65_LH_NAND4ABX3 U9526 ( .A(n7215), .B(n7214), .C(n7213), .D(n7212), .Z(
        n7221) );
  HS65_LH_NAND4ABX3 U9527 ( .A(n7219), .B(n7218), .C(n7217), .D(n7216), .Z(
        n7220) );
  HS65_LH_NOR4ABX2 U9528 ( .A(n7227), .B(n7226), .C(n7225), .D(n7224), .Z(
        n7243) );
  HS65_LH_AOI22X1 U9529 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][23] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][23] ), .D(
        n6957), .Z(n7230) );
  HS65_LH_NOR4ABX2 U9530 ( .A(n7231), .B(n7230), .C(n7229), .D(n7228), .Z(
        n7242) );
  HS65_LH_NAND4ABX3 U9531 ( .A(n7235), .B(n7234), .C(n7233), .D(n7232), .Z(
        n7241) );
  HS65_LH_NAND4ABX3 U9532 ( .A(n7239), .B(n7238), .C(n7237), .D(n7236), .Z(
        n7240) );
  HS65_LH_NOR4ABX2 U9533 ( .A(n7247), .B(n7246), .C(n7245), .D(n7244), .Z(
        n7263) );
  HS65_LH_AOI22X1 U9534 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][6] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][6] ), .D(n6957), .Z(n7250) );
  HS65_LH_NOR4ABX2 U9535 ( .A(n7251), .B(n7250), .C(n7249), .D(n7248), .Z(
        n7262) );
  HS65_LH_NAND4ABX3 U9536 ( .A(n7255), .B(n7254), .C(n7253), .D(n7252), .Z(
        n7261) );
  HS65_LH_NAND4ABX3 U9537 ( .A(n7259), .B(n7258), .C(n7257), .D(n7256), .Z(
        n7260) );
  HS65_LH_AO22X9 U9538 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][29] ), .B(n6364), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][29] ), .D(
        n7266), .Z(n7269) );
  HS65_LH_NOR4ABX2 U9540 ( .A(n7271), .B(n7270), .C(n7269), .D(n7268), .Z(
        n7305) );
  HS65_LH_AO22X9 U9541 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][29] ), .D(
        n7274), .Z(n7279) );
  HS65_LH_AO22X9 U9542 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][29] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][29] ), .D(
        n7276), .Z(n7278) );
  HS65_LH_NOR4ABX2 U9543 ( .A(n7281), .B(n7280), .C(n7279), .D(n7278), .Z(
        n7304) );
  HS65_LH_NAND4ABX3 U9544 ( .A(n7290), .B(n7289), .C(n7288), .D(n7287), .Z(
        n7303) );
  HS65_LH_AO22X9 U9545 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][29] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][29] ), .D(
        n7291), .Z(n7301) );
  HS65_LH_AOI22X1 U9546 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][29] ), .B(n7295), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][29] ), .D(
        n7294), .Z(n7299) );
  HS65_LH_NAND4ABX3 U9547 ( .A(n7301), .B(n7300), .C(n7299), .D(n7298), .Z(
        n7302) );
  HS65_LH_NOR4ABX2 U9548 ( .A(n7305), .B(n7304), .C(n7303), .D(n7302), .Z(
        n8448) );
  HS65_LH_NOR2X2 U9549 ( .A(n8550), .B(n9401), .Z(n8551) );
  HS65_LH_CNIVX3 U9550 ( .A(n7694), .Z(n7772) );
  HS65_LH_NOR4ABX2 U9551 ( .A(n7316), .B(n7315), .C(n7314), .D(n7313), .Z(
        n7342) );
  HS65_LH_AOI22X1 U9552 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][26] ), .B(n7317), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][26] ), .D(
        n6957), .Z(n7323) );
  HS65_LH_NOR4ABX2 U9553 ( .A(n7324), .B(n7323), .C(n7322), .D(n7321), .Z(
        n7341) );
  HS65_LH_NAND4ABX3 U9554 ( .A(n7328), .B(n7327), .C(n7326), .D(n7325), .Z(
        n7340) );
  HS65_LH_NAND4ABX3 U9555 ( .A(n7338), .B(n7337), .C(n7336), .D(n7335), .Z(
        n7339) );
  HS65_LH_NAND2X2 U9556 ( .A(n7343), .B(n7089), .Z(n8146) );
  HS65_LH_NOR4ABX2 U9559 ( .A(n7350), .B(n7349), .C(n7348), .D(n7347), .Z(
        n7366) );
  HS65_LH_NOR4ABX2 U9560 ( .A(n7354), .B(n7353), .C(n7352), .D(n7351), .Z(
        n7365) );
  HS65_LH_NAND4ABX3 U9561 ( .A(n7358), .B(n7357), .C(n7356), .D(n7355), .Z(
        n7364) );
  HS65_LH_NAND4ABX3 U9562 ( .A(n7362), .B(n7361), .C(n7360), .D(n7359), .Z(
        n7363) );
  HS65_LH_NOR4ABX2 U9563 ( .A(n7370), .B(n7369), .C(n7368), .D(n7367), .Z(
        n7386) );
  HS65_LH_NOR4ABX2 U9564 ( .A(n7374), .B(n7373), .C(n7372), .D(n7371), .Z(
        n7385) );
  HS65_LH_NAND4ABX3 U9565 ( .A(n7378), .B(n7377), .C(n7376), .D(n7375), .Z(
        n7384) );
  HS65_LH_NAND4ABX3 U9566 ( .A(n7382), .B(n7381), .C(n7380), .D(n7379), .Z(
        n7383) );
  HS65_LH_NOR4ABX2 U9567 ( .A(n7390), .B(n7389), .C(n7388), .D(n7387), .Z(
        n7406) );
  HS65_LH_NOR4ABX2 U9568 ( .A(n7394), .B(n7393), .C(n7392), .D(n7391), .Z(
        n7405) );
  HS65_LH_NAND4ABX3 U9569 ( .A(n7398), .B(n7397), .C(n7396), .D(n7395), .Z(
        n7404) );
  HS65_LH_NAND4ABX3 U9570 ( .A(n7402), .B(n7401), .C(n7400), .D(n7399), .Z(
        n7403) );
  HS65_LH_NOR4ABX2 U9571 ( .A(n7410), .B(n7409), .C(n7408), .D(n7407), .Z(
        n7427) );
  HS65_LH_NOR4ABX2 U9572 ( .A(n7414), .B(n7413), .C(n7412), .D(n7411), .Z(
        n7426) );
  HS65_LH_NAND4ABX3 U9573 ( .A(n7419), .B(n7418), .C(n7417), .D(n7416), .Z(
        n7425) );
  HS65_LH_NAND4ABX3 U9574 ( .A(n7423), .B(n7422), .C(n7421), .D(n7420), .Z(
        n7424) );
  HS65_LH_NOR4ABX2 U9575 ( .A(n7433), .B(n7432), .C(n7431), .D(n7430), .Z(
        n7451) );
  HS65_LH_NOR4ABX2 U9576 ( .A(n7438), .B(n7437), .C(n7436), .D(n7435), .Z(
        n7450) );
  HS65_LH_NAND4ABX3 U9577 ( .A(n7443), .B(n7442), .C(n7441), .D(n7440), .Z(
        n7449) );
  HS65_LH_NAND4ABX3 U9578 ( .A(n7447), .B(n7446), .C(n7445), .D(n7444), .Z(
        n7448) );
  HS65_LH_NOR4ABX2 U9579 ( .A(n7455), .B(n7454), .C(n7453), .D(n7452), .Z(
        n7471) );
  HS65_LH_NOR4ABX2 U9580 ( .A(n7459), .B(n7458), .C(n7457), .D(n7456), .Z(
        n7470) );
  HS65_LH_NAND4ABX3 U9581 ( .A(n7463), .B(n7462), .C(n7461), .D(n7460), .Z(
        n7469) );
  HS65_LH_NAND4ABX3 U9582 ( .A(n7467), .B(n7466), .C(n7465), .D(n7464), .Z(
        n7468) );
  HS65_LH_AOI22X1 U9583 ( .A(n6739), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][20] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[0][20] ), .D(n6740), 
        .Z(n7474) );
  HS65_LH_NOR4ABX2 U9584 ( .A(n7475), .B(n7474), .C(n7473), .D(n7472), .Z(
        n7491) );
  HS65_LH_NOR4ABX2 U9585 ( .A(n7479), .B(n7478), .C(n7477), .D(n7476), .Z(
        n7490) );
  HS65_LH_NAND4ABX3 U9586 ( .A(n7483), .B(n7482), .C(n7481), .D(n7480), .Z(
        n7489) );
  HS65_LH_NAND4ABX3 U9587 ( .A(n7487), .B(n7486), .C(n7485), .D(n7484), .Z(
        n7488) );
  HS65_LH_NOR4ABX2 U9588 ( .A(n7495), .B(n7494), .C(n7493), .D(n7492), .Z(
        n7511) );
  HS65_LH_NOR4ABX2 U9589 ( .A(n7499), .B(n7498), .C(n7497), .D(n7496), .Z(
        n7510) );
  HS65_LH_NAND4ABX3 U9590 ( .A(n7503), .B(n7502), .C(n7501), .D(n7500), .Z(
        n7509) );
  HS65_LH_NAND4ABX3 U9591 ( .A(n7507), .B(n7506), .C(n7505), .D(n7504), .Z(
        n7508) );
  HS65_LH_NOR4ABX2 U9592 ( .A(n7515), .B(n7514), .C(n7513), .D(n7512), .Z(
        n7537) );
  HS65_LH_NOR4ABX2 U9593 ( .A(n7521), .B(n7520), .C(n7519), .D(n7518), .Z(
        n7536) );
  HS65_LH_NAND4ABX3 U9594 ( .A(n7529), .B(n7528), .C(n7527), .D(n7526), .Z(
        n7535) );
  HS65_LH_NAND4ABX3 U9595 ( .A(n7533), .B(n7532), .C(n7531), .D(n7530), .Z(
        n7534) );
  HS65_LH_NOR4ABX2 U9596 ( .A(n7541), .B(n7540), .C(n7539), .D(n7538), .Z(
        n7557) );
  HS65_LH_NOR4ABX2 U9597 ( .A(n7545), .B(n7544), .C(n7543), .D(n7542), .Z(
        n7556) );
  HS65_LH_NAND4ABX3 U9598 ( .A(n7549), .B(n7548), .C(n7547), .D(n7546), .Z(
        n7555) );
  HS65_LH_NAND4ABX3 U9599 ( .A(n7553), .B(n7552), .C(n7551), .D(n7550), .Z(
        n7554) );
  HS65_LH_NOR4ABX2 U9600 ( .A(n7561), .B(n7560), .C(n7559), .D(n7558), .Z(
        n7577) );
  HS65_LH_NOR4ABX2 U9601 ( .A(n7565), .B(n7564), .C(n7563), .D(n7562), .Z(
        n7576) );
  HS65_LH_NAND4ABX3 U9602 ( .A(n7569), .B(n7568), .C(n7567), .D(n7566), .Z(
        n7575) );
  HS65_LH_NAND4ABX3 U9603 ( .A(n7573), .B(n7572), .C(n7571), .D(n7570), .Z(
        n7574) );
  HS65_LH_NOR4ABX2 U9604 ( .A(n7584), .B(n7583), .C(n7582), .D(n7581), .Z(
        n7612) );
  HS65_LH_NOR4ABX2 U9605 ( .A(n7591), .B(n7590), .C(n7589), .D(n7588), .Z(
        n7611) );
  HS65_LH_NAND4ABX3 U9606 ( .A(n7598), .B(n7597), .C(n7596), .D(n7595), .Z(
        n7610) );
  HS65_LH_NAND4ABX3 U9607 ( .A(n7608), .B(n7607), .C(n7606), .D(n7605), .Z(
        n7609) );
  HS65_LH_NOR2X2 U9608 ( .A(\u_DataPath/u_idexreg/N3 ), .B(n7617), .Z(
        \u_DataPath/u_execute/EXALU/N810 ) );
  HS65_LH_IVX2 U9609 ( .A(n7618), .Z(n8138) );
  HS65_LH_IVX2 U9610 ( .A(n7619), .Z(n8142) );
  HS65_LH_NOR2AX3 U9611 ( .A(n9076), .B(n2847), .Z(n7733) );
  HS65_LH_NAND2X2 U9612 ( .A(n7733), .B(n9031), .Z(n8149) );
  HS65_LH_NOR2X2 U9613 ( .A(n2851), .B(n7621), .Z(n7625) );
  HS65_LH_NOR2X2 U9614 ( .A(n7622), .B(n2840), .Z(n7624) );
  HS65_LH_MUXI21X2 U9615 ( .D0(n7625), .D1(n7624), .S0(n7623), .Z(n7635) );
  HS65_LH_NAND2X2 U9616 ( .A(n7626), .B(n2840), .Z(n7629) );
  HS65_LH_NOR2X2 U9617 ( .A(n7626), .B(n2840), .Z(n7628) );
  HS65_LH_MUX21I1X3 U9618 ( .D0(n7629), .D1(n7628), .S0(n7627), .Z(n7630) );
  HS65_LH_NAND2X2 U9619 ( .A(n7631), .B(n7630), .Z(n7633) );
  HS65_LH_CBI4I6X2 U9620 ( .A(n7635), .B(n7634), .C(n7633), .D(
        \u_DataPath/u_idexreg/N3 ), .Z(\u_DataPath/u_execute/EXALU/N811 ) );
  HS65_LH_CNIVX3 U9621 ( .A(\u_DataPath/jaddr_i [19]), .Z(n8042) );
  HS65_LH_IVX2 U9622 ( .A(n8716), .Z(n8490) );
  HS65_LH_IVX2 U9624 ( .A(Data_out_fromRAM[18]), .Z(n8454) );
  HS65_LH_IVX2 U9625 ( .A(Data_out_fromRAM[19]), .Z(n8324) );
  HS65_LH_IVX2 U9626 ( .A(Data_out_fromRAM[22]), .Z(n8351) );
  HS65_LH_IVX2 U9627 ( .A(Data_out_fromRAM[16]), .Z(n8356) );
  HS65_LH_IVX2 U9628 ( .A(Data_out_fromRAM[17]), .Z(n8406) );
  HS65_LH_NOR2X6 U9631 ( .A(n7648), .B(n7676), .Z(n7649) );
  HS65_LH_CNIVX3 U9632 ( .A(n7652), .Z(n7654) );
  HS65_LH_NOR2X2 U9635 ( .A(opcode_i[1]), .B(opcode_i[3]), .Z(n7696) );
  HS65_LH_CNIVX3 U9636 ( .A(n8086), .Z(n7702) );
  HS65_LH_NOR3X1 U9637 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .B(
        \u_DataPath/immediate_ext_dec_i [3]), .C(n8092), .Z(n7699) );
  HS65_LH_NAND2X2 U9638 ( .A(n8076), .B(n7699), .Z(n7701) );
  HS65_LH_CNIVX3 U9639 ( .A(n8076), .Z(n7703) );
  HS65_LH_NAND4ABX3 U9640 ( .A(opcode_i[3]), .B(n9082), .C(n7735), .D(n7778), 
        .Z(n8049) );
  HS65_LH_NOR3X1 U9641 ( .A(\u_DataPath/immediate_ext_dec_i [2]), .B(
        \u_DataPath/immediate_ext_dec_i [3]), .C(
        \u_DataPath/immediate_ext_dec_i [10]), .Z(n7737) );
  HS65_LH_NOR2X2 U9642 ( .A(\u_DataPath/immediate_ext_dec_i [8]), .B(
        \u_DataPath/immediate_ext_dec_i [9]), .Z(n7736) );
  HS65_LH_NAND4ABX3 U9643 ( .A(\u_DataPath/immediate_ext_dec_i [6]), .B(
        \u_DataPath/immediate_ext_dec_i [7]), .C(n7737), .D(n7736), .Z(n8073)
         );
  HS65_LH_NAND4ABX3 U9644 ( .A(n7763), .B(n7740), .C(n7739), .D(n8083), .Z(
        n8057) );
  HS65_LH_NAND4ABX3 U9646 ( .A(n8123), .B(n8122), .C(n8121), .D(n8120), .Z(
        n7760) );
  HS65_LH_AOI21X2 U9647 ( .A(n7772), .B(n7777), .C(n7763), .Z(n8100) );
  HS65_LH_AOI21X2 U9648 ( .A(n7773), .B(n7772), .C(n7771), .Z(n7774) );
  HS65_LH_AOI222X2 U9649 ( .A(n7779), .B(opcode_i[1]), .C(n7778), .D(n7777), 
        .E(n9084), .F(n7776), .Z(n8081) );
  HS65_LH_HA1X4 U9650 ( .A0(n2908), .B0(n9204), .CO(n7801), .S0(
        \u_DataPath/u_execute/link_value_i [29]) );
  HS65_LH_HA1X4 U9651 ( .A0(n7801), .B0(n9203), .CO(n7800), .S0(
        \u_DataPath/u_execute/link_value_i [30]) );
  HS65_LH_NOR2X2 U9652 ( .A(n8840), .B(n7802), .Z(n7803) );
  HS65_LH_AND2X4 U9653 ( .A(n2896), .B(n7803), .Z(n7864) );
  HS65_LL_OAI21X18 U9655 ( .A(n3009), .B(n8141), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N148 ) );
  HS65_LL_OAI21X18 U9656 ( .A(n3010), .B(n8141), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N153 ) );
  HS65_LL_OAI21X12 U9657 ( .A(n8141), .B(n2773), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N149 ) );
  HS65_LL_OAI21X12 U9658 ( .A(n8150), .B(n8145), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N133 ) );
  HS65_LL_OAI21X12 U9659 ( .A(n8150), .B(n3012), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N134 ) );
  HS65_LL_OAI21X12 U9660 ( .A(n8141), .B(n3012), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N150 ) );
  HS65_LL_OAI21X12 U9661 ( .A(n8140), .B(n3012), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N142 ) );
  HS65_LH_NOR2X2 U9662 ( .A(rst), .B(n8160), .Z(
        \u_DataPath/u_decode_unit/hdu_0/current_state [1]) );
  HS65_LH_BFX18 U9663 ( .A(n8443), .Z(n7899) );
  HS65_LH_BFX18 U9664 ( .A(n8443), .Z(n7900) );
  HS65_LH_NAND3X3 U9665 ( .A(n8142), .B(n8143), .C(n8139), .Z(n8141) );
  HS65_LH_NAND3X2 U9666 ( .A(n9075), .B(n8138), .C(n8143), .Z(n8140) );
  HS65_LH_AND2X4 U9667 ( .A(n2733), .B(\u_DataPath/toPC2_i [24]), .Z(
        \u_DataPath/branch_target_i [24]) );
  HS65_LH_NOR4ABX2 U9668 ( .A(n8566), .B(n8565), .C(n8564), .D(n7878), .Z(
        \u_DataPath/mem_writedata_out_i [29]) );
  HS65_LH_NOR4ABX2 U9669 ( .A(n8566), .B(n8560), .C(n8559), .D(n8558), .Z(
        \u_DataPath/mem_writedata_out_i [27]) );
  HS65_LH_NOR4ABX2 U9670 ( .A(n8566), .B(n8540), .C(n8539), .D(n8538), .Z(
        \u_DataPath/mem_writedata_out_i [20]) );
  HS65_LH_NOR4ABX2 U9671 ( .A(n8566), .B(n8543), .C(n8542), .D(n8541), .Z(
        \u_DataPath/mem_writedata_out_i [21]) );
  HS65_LH_AND2X4 U9674 ( .A(n2733), .B(\u_DataPath/toPC2_i [15]), .Z(
        \u_DataPath/branch_target_i [15]) );
  HS65_LH_AO222X4 U9675 ( .A(n7895), .B(\u_DataPath/pc_4_i [12]), .C(n7892), 
        .D(n9412), .E(n8917), .F(n7888), .Z(n8660) );
  HS65_LH_AO222X4 U9676 ( .A(n7895), .B(\u_DataPath/pc_4_i [14]), .C(n7892), 
        .D(\u_DataPath/jump_address_i [14]), .E(n9198), .F(n7888), .Z(n8658)
         );
  HS65_LH_AO222X4 U9677 ( .A(n7895), .B(\u_DataPath/pc_4_i [18]), .C(n7892), 
        .D(n9411), .E(n8927), .F(n7887), .Z(n8654) );
  HS65_LH_AO222X4 U9678 ( .A(n7895), .B(\u_DataPath/pc_4_i [19]), .C(n7892), 
        .D(\u_DataPath/jump_address_i [19]), .E(n8925), .F(n7887), .Z(n8653)
         );
  HS65_LH_NOR3AX4 U9679 ( .A(n8755), .B(rst), .C(\u_DataPath/cw_to_ex_i [15]), 
        .Z(n8450) );
  HS65_LH_NOR4ABX2 U9680 ( .A(n8566), .B(n8502), .C(n8501), .D(n8500), .Z(
        \u_DataPath/mem_writedata_out_i [7]) );
  HS65_LH_NOR4ABX2 U9681 ( .A(n8566), .B(n8486), .C(n7864), .D(n8485), .Z(
        \u_DataPath/mem_writedata_out_i [1]) );
  HS65_LH_NOR4ABX2 U9682 ( .A(n8566), .B(n8499), .C(n8498), .D(n8497), .Z(
        \u_DataPath/mem_writedata_out_i [6]) );
  HS65_LH_NOR4ABX2 U9683 ( .A(n8518), .B(n8517), .C(n8516), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [13]) );
  HS65_LH_NOR4ABX2 U9684 ( .A(n8509), .B(n8508), .C(n8507), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [10]) );
  HS65_LH_NOR4ABX2 U9685 ( .A(n8530), .B(n8529), .C(n8528), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [17]) );
  HS65_LH_NOR4ABX2 U9686 ( .A(n8521), .B(n8520), .C(n8519), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [14]) );
  HS65_LH_NOR4ABX2 U9687 ( .A(n8527), .B(n8526), .C(n8525), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [16]) );
  HS65_LH_NOR4ABX2 U9688 ( .A(n8533), .B(n8532), .C(n8531), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [18]) );
  HS65_LH_NOR4ABX2 U9689 ( .A(n8549), .B(n8548), .C(n8547), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [23]) );
  HS65_LH_NOR4ABX2 U9690 ( .A(n8512), .B(n8511), .C(n8510), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [11]) );
  HS65_LH_NOR4ABX2 U9691 ( .A(n8524), .B(n8523), .C(n8522), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [15]) );
  HS65_LH_NOR4ABX2 U9692 ( .A(n8557), .B(n8556), .C(n8555), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [26]) );
  HS65_LH_NOR4ABX2 U9693 ( .A(n8553), .B(n8552), .C(rst), .D(n8551), .Z(
        \u_DataPath/mem_writedata_out_i [24]) );
  HS65_LH_NOR4ABX2 U9694 ( .A(n8496), .B(n8495), .C(n7863), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [5]) );
  HS65_LH_NOR4ABX2 U9695 ( .A(n8515), .B(n8514), .C(n8513), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [12]) );
  HS65_LH_NOR4ABX2 U9696 ( .A(n8569), .B(n8568), .C(n8567), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [30]) );
  HS65_LH_NOR4ABX2 U9697 ( .A(n8572), .B(n8571), .C(n8570), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [31]) );
  HS65_LH_NOR4ABX2 U9698 ( .A(n8546), .B(n8545), .C(n8544), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [22]) );
  HS65_LH_AND2X4 U9699 ( .A(n2733), .B(\u_DataPath/toPC2_i [22]), .Z(
        \u_DataPath/branch_target_i [22]) );
  HS65_LH_AND2X4 U9700 ( .A(n2733), .B(\u_DataPath/toPC2_i [17]), .Z(
        \u_DataPath/branch_target_i [17]) );
  HS65_LH_AND2X4 U9701 ( .A(n2733), .B(\u_DataPath/toPC2_i [18]), .Z(
        \u_DataPath/branch_target_i [18]) );
  HS65_LH_AND2X4 U9702 ( .A(n2733), .B(\u_DataPath/toPC2_i [20]), .Z(
        \u_DataPath/branch_target_i [20]) );
  HS65_LH_AND2X4 U9703 ( .A(n2733), .B(\u_DataPath/toPC2_i [19]), .Z(
        \u_DataPath/branch_target_i [19]) );
  HS65_LH_NOR2X2 U9704 ( .A(n8262), .B(rst), .Z(n8143) );
  HS65_LH_BFX4 U9705 ( .A(n8609), .Z(n8004) );
  HS65_LH_BFX4 U9706 ( .A(n8607), .Z(n7995) );
  HS65_LH_BFX4 U9707 ( .A(n8599), .Z(n7968) );
  HS65_LH_BFX4 U9708 ( .A(n8593), .Z(n7950) );
  HS65_LH_BFX4 U9709 ( .A(n8595), .Z(n7956) );
  HS65_LH_BFX4 U9710 ( .A(n8610), .Z(n8007) );
  HS65_LH_BFX4 U9711 ( .A(n8598), .Z(n7965) );
  HS65_LH_BFX4 U9712 ( .A(n8616), .Z(n8022) );
  HS65_LH_BFX4 U9713 ( .A(n8606), .Z(n7992) );
  HS65_LH_BFX4 U9714 ( .A(n8612), .Z(n8013) );
  HS65_LH_BFX4 U9715 ( .A(n8603), .Z(n7983) );
  HS65_LH_BFX4 U9716 ( .A(n8601), .Z(n7977) );
  HS65_LH_BFX4 U9717 ( .A(n8622), .Z(n8031) );
  HS65_LH_BFX4 U9718 ( .A(n8588), .Z(n7938) );
  HS65_LH_BFX4 U9719 ( .A(n8596), .Z(n7959) );
  HS65_LH_BFX4 U9720 ( .A(n8594), .Z(n7953) );
  HS65_LH_BFX4 U9721 ( .A(n8604), .Z(n7986) );
  HS65_LH_BFX4 U9722 ( .A(n8620), .Z(n8028) );
  HS65_LH_BFX4 U9723 ( .A(n8602), .Z(n7980) );
  HS65_LH_BFX4 U9724 ( .A(n8613), .Z(n8016) );
  HS65_LH_BFX4 U9725 ( .A(n8618), .Z(n8025) );
  HS65_LH_BFX4 U9726 ( .A(n8611), .Z(n8011) );
  HS65_LH_BFX4 U9727 ( .A(n8611), .Z(n8012) );
  HS65_LH_BFX4 U9728 ( .A(n8587), .Z(n7935) );
  HS65_LH_CNIVX3 U9729 ( .A(n8608), .Z(n8003) );
  HS65_LH_BFX4 U9730 ( .A(n8585), .Z(n7928) );
  HS65_LH_BFX4 U9731 ( .A(n8605), .Z(n7991) );
  HS65_LH_BFX4 U9732 ( .A(n8589), .Z(n7943) );
  HS65_LH_BFX4 U9733 ( .A(n8597), .Z(n7964) );
  HS65_LH_BFX4 U9734 ( .A(n8614), .Z(n8021) );
  HS65_LH_BFX4 U9735 ( .A(n8609), .Z(n8006) );
  HS65_LH_BFX4 U9736 ( .A(n8607), .Z(n7997) );
  HS65_LH_BFX4 U9737 ( .A(n8599), .Z(n7970) );
  HS65_LH_BFX4 U9738 ( .A(n8614), .Z(n8019) );
  HS65_LH_BFX4 U9739 ( .A(n8597), .Z(n7962) );
  HS65_LH_BFX4 U9740 ( .A(n8589), .Z(n7941) );
  HS65_LH_CNIVX3 U9741 ( .A(n8600), .Z(n7976) );
  HS65_LH_BFX4 U9742 ( .A(n8605), .Z(n7989) );
  HS65_LH_BFX4 U9743 ( .A(n8585), .Z(n7926) );
  HS65_LH_BFX4 U9744 ( .A(n8587), .Z(n7936) );
  HS65_LH_CNIVX3 U9745 ( .A(n8608), .Z(n8002) );
  HS65_LH_BFX4 U9746 ( .A(n8618), .Z(n8026) );
  HS65_LH_BFX4 U9747 ( .A(n8613), .Z(n8017) );
  HS65_LH_BFX4 U9748 ( .A(n8602), .Z(n7981) );
  HS65_LH_BFX4 U9749 ( .A(n8620), .Z(n8029) );
  HS65_LH_BFX4 U9750 ( .A(n8604), .Z(n7987) );
  HS65_LH_BFX4 U9751 ( .A(n8594), .Z(n7954) );
  HS65_LH_BFX4 U9752 ( .A(n8596), .Z(n7960) );
  HS65_LH_BFX4 U9753 ( .A(n8588), .Z(n7939) );
  HS65_LH_BFX4 U9754 ( .A(n8622), .Z(n8032) );
  HS65_LH_BFX4 U9755 ( .A(n8601), .Z(n7978) );
  HS65_LH_BFX4 U9756 ( .A(n8603), .Z(n7984) );
  HS65_LH_BFX4 U9757 ( .A(n8612), .Z(n8014) );
  HS65_LH_BFX4 U9758 ( .A(n8606), .Z(n7993) );
  HS65_LH_BFX4 U9759 ( .A(n8616), .Z(n8023) );
  HS65_LH_BFX4 U9760 ( .A(n8598), .Z(n7966) );
  HS65_LH_BFX4 U9761 ( .A(n8610), .Z(n8008) );
  HS65_LH_BFX4 U9762 ( .A(n8595), .Z(n7957) );
  HS65_LH_BFX4 U9763 ( .A(n8593), .Z(n7951) );
  HS65_LH_BFX4 U9764 ( .A(n8599), .Z(n7969) );
  HS65_LH_CNIVX3 U9765 ( .A(n8293), .Z(n8599) );
  HS65_LH_BFX4 U9766 ( .A(n8611), .Z(n8010) );
  HS65_LH_CNIVX3 U9767 ( .A(n8397), .Z(n8611) );
  HS65_LH_BFX4 U9768 ( .A(n8607), .Z(n7996) );
  HS65_LH_CNIVX3 U9769 ( .A(n8362), .Z(n8607) );
  HS65_LH_BFX4 U9770 ( .A(n8609), .Z(n8005) );
  HS65_LH_CNIVX3 U9771 ( .A(n8321), .Z(n8609) );
  HS65_LH_CNIVX3 U9772 ( .A(n8591), .Z(n7948) );
  HS65_LH_BFX4 U9773 ( .A(n8614), .Z(n8020) );
  HS65_LH_CNIVX3 U9774 ( .A(n8434), .Z(n8614) );
  HS65_LH_BFX4 U9775 ( .A(n8597), .Z(n7963) );
  HS65_LH_CNIVX3 U9776 ( .A(n8326), .Z(n8597) );
  HS65_LH_BFX4 U9777 ( .A(n8589), .Z(n7942) );
  HS65_LH_CNIVX3 U9778 ( .A(n8348), .Z(n8589) );
  HS65_LH_CNIVX3 U9779 ( .A(n8600), .Z(n7975) );
  HS65_LH_BFX4 U9780 ( .A(n8605), .Z(n7990) );
  HS65_LH_CNIVX3 U9781 ( .A(n8404), .Z(n8605) );
  HS65_LH_BFX4 U9782 ( .A(n8585), .Z(n7927) );
  HS65_LH_CNIVX3 U9783 ( .A(n8378), .Z(n8585) );
  HS65_LH_BFX4 U9784 ( .A(n8587), .Z(n7937) );
  HS65_LH_CNIVX3 U9785 ( .A(n8422), .Z(n8587) );
  HS65_LH_BFX4 U9786 ( .A(n8618), .Z(n8027) );
  HS65_LH_CNIVX3 U9787 ( .A(n8168), .Z(n8618) );
  HS65_LH_CNIVX3 U9788 ( .A(n8591), .Z(n7949) );
  HS65_LH_BFX4 U9789 ( .A(n8613), .Z(n8018) );
  HS65_LH_CNIVX3 U9790 ( .A(n8314), .Z(n8613) );
  HS65_LH_BFX4 U9791 ( .A(n8593), .Z(n7952) );
  HS65_LH_CNIVX3 U9792 ( .A(n8304), .Z(n8593) );
  HS65_LH_BFX4 U9793 ( .A(n8595), .Z(n7958) );
  HS65_LH_CNIVX3 U9794 ( .A(n8343), .Z(n8595) );
  HS65_LH_BFX4 U9795 ( .A(n8610), .Z(n8009) );
  HS65_LH_CNIVX3 U9796 ( .A(n8449), .Z(n8610) );
  HS65_LH_BFX4 U9797 ( .A(n8598), .Z(n7967) );
  HS65_LH_CNIVX3 U9798 ( .A(n8367), .Z(n8598) );
  HS65_LH_BFX4 U9799 ( .A(n8602), .Z(n7982) );
  HS65_LH_CNIVX3 U9800 ( .A(n8457), .Z(n8602) );
  HS65_LH_BFX4 U9801 ( .A(n8616), .Z(n8024) );
  HS65_LH_CNIVX3 U9802 ( .A(n8415), .Z(n8616) );
  HS65_LH_BFX4 U9803 ( .A(n8606), .Z(n7994) );
  HS65_LH_CNIVX3 U9804 ( .A(n8330), .Z(n8606) );
  HS65_LH_BFX4 U9805 ( .A(n8612), .Z(n8015) );
  HS65_LH_CNIVX3 U9806 ( .A(n8337), .Z(n8612) );
  HS65_LH_BFX4 U9807 ( .A(n8603), .Z(n7985) );
  HS65_LH_CNIVX3 U9808 ( .A(n8372), .Z(n8603) );
  HS65_LH_BFX4 U9809 ( .A(n8596), .Z(n7961) );
  HS65_LH_CNIVX3 U9810 ( .A(n8412), .Z(n8596) );
  HS65_LH_BFX4 U9811 ( .A(n8622), .Z(n8033) );
  HS65_LH_CNIVX3 U9812 ( .A(n8431), .Z(n8622) );
  HS65_LH_BFX4 U9813 ( .A(n8604), .Z(n7988) );
  HS65_LH_CNIVX3 U9814 ( .A(n8408), .Z(n8604) );
  HS65_LH_BFX4 U9815 ( .A(n8620), .Z(n8030) );
  HS65_LH_CNIVX3 U9816 ( .A(n8444), .Z(n8620) );
  HS65_LH_BFX4 U9817 ( .A(n8594), .Z(n7955) );
  HS65_LH_CNIVX3 U9818 ( .A(n8358), .Z(n8594) );
  HS65_LH_BFX4 U9819 ( .A(n8588), .Z(n7940) );
  HS65_LH_CNIVX3 U9820 ( .A(n8275), .Z(n8588) );
  HS65_LH_BFX4 U9821 ( .A(n8601), .Z(n7979) );
  HS65_LH_CNIVX3 U9822 ( .A(n8353), .Z(n8601) );
  HS65_LH_AND2X4 U9823 ( .A(n2733), .B(\u_DataPath/toPC2_i [1]), .Z(
        \u_DataPath/branch_target_i [1]) );
  HS65_LH_NOR4ABX2 U9824 ( .A(n8506), .B(n8505), .C(n8504), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [9]) );
  HS65_LH_AND2X4 U9825 ( .A(n2733), .B(\u_DataPath/toPC2_i [2]), .Z(
        \u_DataPath/branch_target_i [2]) );
  HS65_LH_NOR4ABX2 U9826 ( .A(n8492), .B(n8491), .C(n3312), .D(rst), .Z(
        \u_DataPath/mem_writedata_out_i [3]) );
  HS65_LH_NOR2X2 U9827 ( .A(rst), .B(n8034), .Z(
        \u_DataPath/u_decode_unit/hdu_0/current_state [0]) );
  HS65_LH_AND2X4 U9828 ( .A(n2733), .B(\u_DataPath/toPC2_i [5]), .Z(
        \u_DataPath/branch_target_i [5]) );
  HS65_LH_AND2X4 U9829 ( .A(n2733), .B(\u_DataPath/toPC2_i [6]), .Z(
        \u_DataPath/branch_target_i [6]) );
  HS65_LH_AND2X4 U9830 ( .A(n2733), .B(\u_DataPath/toPC2_i [8]), .Z(
        \u_DataPath/branch_target_i [8]) );
  HS65_LH_AND2X4 U9831 ( .A(n2733), .B(\u_DataPath/toPC2_i [13]), .Z(
        \u_DataPath/branch_target_i [13]) );
  HS65_LH_AND2X4 U9832 ( .A(n2733), .B(\u_DataPath/toPC2_i [11]), .Z(
        \u_DataPath/branch_target_i [11]) );
  HS65_LH_AND2X4 U9833 ( .A(n2733), .B(\u_DataPath/toPC2_i [12]), .Z(
        \u_DataPath/branch_target_i [12]) );
  HS65_LH_OAI12X6 U9834 ( .A(n8140), .B(n8149), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N144 ) );
  HS65_LH_OAI12X6 U9835 ( .A(n8141), .B(n8149), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N152 ) );
  HS65_LH_OAI12X6 U9836 ( .A(n8144), .B(n8150), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N138 ) );
  HS65_LH_OAI12X6 U9837 ( .A(n8144), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N130 ) );
  HS65_LH_OAI12X6 U9838 ( .A(n8146), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N131 ) );
  HS65_LH_OAI12X6 U9839 ( .A(n8140), .B(n8144), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N146 ) );
  HS65_LH_OAI12X6 U9840 ( .A(n8149), .B(n8150), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N136 ) );
  HS65_LH_OAI12X6 U9841 ( .A(n8144), .B(n8141), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N154 ) );
  HS65_LH_OAI12X6 U9842 ( .A(n8140), .B(n8146), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N147 ) );
  HS65_LH_OAI12X6 U9843 ( .A(n8146), .B(n8150), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N139 ) );
  HS65_LH_NAND3X5 U9844 ( .A(n8960), .B(n8142), .C(n8143), .Z(n8150) );
  HS65_LH_OAI12X6 U9845 ( .A(n8149), .B(n8148), .C(n2733), .Z(
        \u_DataPath/u_decode_unit/reg_file0/N128 ) );
  HS65_LH_CNIVX3 U9846 ( .A(n7934), .Z(n7929) );
  HS65_LH_CNIVX3 U9847 ( .A(n8586), .Z(n7934) );
  HS65_LH_CNIVX3 U9848 ( .A(n8003), .Z(n7998) );
  HS65_LH_CNIVX3 U9849 ( .A(n7974), .Z(n7973) );
  HS65_LH_CNIVX3 U9850 ( .A(n7947), .Z(n7946) );
  HS65_LH_CNIVX3 U9851 ( .A(n7976), .Z(n7971) );
  HS65_LH_CNIVX3 U9852 ( .A(n8002), .Z(n7999) );
  HS65_LH_CNIVX3 U9853 ( .A(n7933), .Z(n7930) );
  HS65_LH_CNIVX3 U9854 ( .A(n8586), .Z(n7933) );
  HS65_LH_CNIVX3 U9855 ( .A(n7948), .Z(n7945) );
  HS65_LH_CNIVX3 U9856 ( .A(n7975), .Z(n7972) );
  HS65_LH_CNIVX3 U9857 ( .A(n8001), .Z(n8000) );
  HS65_LH_CNIVX3 U9858 ( .A(n7949), .Z(n7944) );
  HS65_LH_CNIVX3 U9859 ( .A(n7932), .Z(n7931) );
  HS65_LH_CNIVX3 U9860 ( .A(n8423), .Z(\u_DataPath/u_execute/psw_status_i [1])
         );
  HS65_LH_CNIVX3 U9864 ( .A(n8228), .Z(\u_DataPath/pc_4_to_ex_i [2]) );
  HS65_LH_CNIVX3 U9865 ( .A(n8230), .Z(\u_DataPath/u_execute/link_value_i [0])
         );
  HS65_LH_CNIVX3 U9866 ( .A(n8113), .Z(\u_DataPath/cw_tomem_i [5]) );
  HS65_LH_CNIVX3 U9867 ( .A(n8109), .Z(\u_DataPath/cw_tomem_i [4]) );
  HS65_LH_CNIVX3 U9868 ( .A(n8061), .Z(\u_DataPath/reg_write_i ) );
  HS65_LH_CNIVX3 U9869 ( .A(n8263), .Z(\u_DataPath/cw_memwb_i [1]) );
  HS65_LH_CNIVX3 U9870 ( .A(n8579), .Z(n8494) );
  HS65_LL_OAI22X1 U9871 ( .A(n7096), .B(n8431), .C(n7901), .D(n8392), .Z(
        \u_DataPath/data_read_ex_2_i [4]) );
  HS65_LL_OAI22X1 U9872 ( .A(n7096), .B(n8404), .C(n7901), .D(n8388), .Z(
        \u_DataPath/data_read_ex_2_i [14]) );
  HS65_LL_OAI22X1 U9873 ( .A(n7096), .B(n8434), .C(n7901), .D(n8433), .Z(
        \u_DataPath/data_read_ex_2_i [3]) );
  HS65_LH_NAND2X7 U9875 ( .A(opcode_i[5]), .B(n8045), .Z(n8053) );
  HS65_LL_OAI22X1 U9876 ( .A(n7096), .B(n8397), .C(n7900), .D(n8379), .Z(
        \u_DataPath/data_read_ex_2_i [30]) );
  HS65_LL_OAI22X1 U9877 ( .A(n7902), .B(n8001), .C(n7899), .D(n8155), .Z(
        \u_DataPath/data_read_ex_2_i [0]) );
  HS65_LL_OAI22X1 U9878 ( .A(n7096), .B(n8378), .C(n7900), .D(n8373), .Z(
        \u_DataPath/data_read_ex_2_i [27]) );
  HS65_LL_OAI22X1 U9879 ( .A(n7096), .B(n8412), .C(n7901), .D(n8384), .Z(
        \u_DataPath/data_read_ex_2_i [20]) );
  HS65_LL_OAI22X1 U9880 ( .A(n7096), .B(n7932), .C(n7901), .D(n8382), .Z(
        \u_DataPath/data_read_ex_2_i [28]) );
  HS65_LL_OAI22X1 U9881 ( .A(n7096), .B(n8449), .C(n7901), .D(n8381), .Z(
        \u_DataPath/data_read_ex_2_i [29]) );
  HS65_LL_OAI22X1 U9882 ( .A(n7096), .B(n8358), .C(n7900), .D(n8354), .Z(
        \u_DataPath/data_read_ex_2_i [16]) );
  HS65_LL_OAI22X1 U9883 ( .A(n7096), .B(n8372), .C(n7900), .D(n8368), .Z(
        \u_DataPath/data_read_ex_2_i [24]) );
  HS65_LL_OAI22X1 U9884 ( .A(n7096), .B(n8367), .C(n7900), .D(n8363), .Z(
        \u_DataPath/data_read_ex_2_i [21]) );
  HS65_LH_OAI211X3 U9885 ( .A(n8696), .B(n9012), .C(n8885), .D(n8079), .Z(
        \u_DataPath/cw_to_ex_i [1]) );
  HS65_LL_OAI22X1 U9888 ( .A(n7096), .B(n8444), .C(n7901), .D(n8442), .Z(
        \u_DataPath/data_read_ex_2_i [2]) );
  HS65_LH_NOR2AX3 U9889 ( .A(n9233), .B(rst), .Z(n8286) );
  HS65_LH_IVX9 U9890 ( .A(n8480), .Z(n7873) );
  HS65_LH_NOR2AX3 U9891 ( .A(\u_DataPath/cw_exmem_i [3]), .B(rst), .Z(
        \u_DataPath/cw_tomem_i [3]) );
  HS65_LH_NOR2AX3 U9892 ( .A(\u_DataPath/dataOut_exe_i [31]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [31]) );
  HS65_LH_NOR2AX3 U9893 ( .A(\u_DataPath/dataOut_exe_i [17]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [17]) );
  HS65_LH_NOR2AX3 U9894 ( .A(\u_DataPath/dataOut_exe_i [16]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [16]) );
  HS65_LH_NOR2AX3 U9895 ( .A(\u_DataPath/dataOut_exe_i [22]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [22]) );
  HS65_LH_NOR2AX3 U9896 ( .A(\u_DataPath/dataOut_exe_i [28]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [28]) );
  HS65_LH_NOR2AX3 U9897 ( .A(\u_DataPath/dataOut_exe_i [9]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [9]) );
  HS65_LH_NOR2AX3 U9898 ( .A(\u_DataPath/dataOut_exe_i [7]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [7]) );
  HS65_LH_NOR2AX3 U9899 ( .A(\u_DataPath/dataOut_exe_i [3]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [3]) );
  HS65_LH_NOR2AX3 U9900 ( .A(\u_DataPath/dataOut_exe_i [29]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [29]) );
  HS65_LH_NOR2AX3 U9901 ( .A(\u_DataPath/dataOut_exe_i [14]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [14]) );
  HS65_LH_NOR2AX3 U9902 ( .A(\u_DataPath/immediate_ext_dec_i [4]), .B(rst), 
        .Z(\u_DataPath/immediate_ext_ex_i [4]) );
  HS65_LH_NOR2X6 U9903 ( .A(n8166), .B(rst), .Z(n8626) );
  HS65_LH_AND2X4 U9904 ( .A(n9068), .B(n8634), .Z(\u_DataPath/cw_to_ex_i [20])
         );
  HS65_LH_MUXI21X2 U9905 ( .D0(n9084), .D1(iram_data[26]), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(n8043) );
  HS65_LH_MUXI21X2 U9906 ( .D0(n9082), .D1(iram_data[28]), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(n8036) );
  HS65_LH_MUXI21X2 U9907 ( .D0(n9068), .D1(iram_data[30]), .S0(
        \u_DataPath/u_fetch/pc1/N3 ), .Z(n8035) );
  HS65_LH_NOR2AX3 U9908 ( .A(\u_DataPath/dataOut_exe_i [15]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [15]) );
  HS65_LH_NOR2AX3 U9909 ( .A(\u_DataPath/dataOut_exe_i [6]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [6]) );
  HS65_LH_NOR2AX3 U9910 ( .A(\u_DataPath/dataOut_exe_i [5]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [5]) );
  HS65_LH_NOR2AX3 U9911 ( .A(\u_DataPath/dataOut_exe_i [23]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [23]) );
  HS65_LH_NOR2AX3 U9912 ( .A(\u_DataPath/dataOut_exe_i [30]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [30]) );
  HS65_LH_NOR2AX3 U9913 ( .A(\u_DataPath/dataOut_exe_i [8]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [8]) );
  HS65_LH_NOR2AX3 U9914 ( .A(\u_DataPath/dataOut_exe_i [26]), .B(rst), .Z(
        \u_DataPath/u_memwbreg/N64 ) );
  HS65_LH_NOR2AX3 U9915 ( .A(\u_DataPath/dataOut_exe_i [24]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [24]) );
  HS65_LH_NOR2AX3 U9916 ( .A(\u_DataPath/dataOut_exe_i [2]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [2]) );
  HS65_LH_NOR2AX3 U9917 ( .A(\u_DataPath/dataOut_exe_i [19]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [19]) );
  HS65_LH_NOR2AX3 U9918 ( .A(\u_DataPath/dataOut_exe_i [18]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [18]) );
  HS65_LH_NOR2AX3 U9919 ( .A(\u_DataPath/dataOut_exe_i [12]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [12]) );
  HS65_LH_NOR2AX3 U9920 ( .A(\u_DataPath/dataOut_exe_i [25]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [25]) );
  HS65_LH_NOR2AX3 U9921 ( .A(\u_DataPath/dataOut_exe_i [13]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [13]) );
  HS65_LH_NOR2AX3 U9922 ( .A(\u_DataPath/dataOut_exe_i [11]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [11]) );
  HS65_LH_NOR2AX3 U9923 ( .A(\u_DataPath/dataOut_exe_i [21]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [21]) );
  HS65_LH_NOR2AX3 U9924 ( .A(\u_DataPath/dataOut_exe_i [27]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [27]) );
  HS65_LH_NOR2AX3 U9925 ( .A(\u_DataPath/dataOut_exe_i [20]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [20]) );
  HS65_LH_NOR2AX3 U9926 ( .A(\u_DataPath/dataOut_exe_i [10]), .B(rst), .Z(
        \u_DataPath/from_alu_data_out_i [10]) );
  HS65_LH_AO22X4 U9927 ( .A(n8580), .B(n8425), .C(n8621), .D(n8573), .Z(
        \u_DataPath/u_execute/psw_status_i [0]) );
  HS65_LH_AO222X4 U9928 ( .A(n7894), .B(n8691), .C(n7891), .D(
        \u_DataPath/jump_address_i [0]), .E(n9250), .F(n7889), .Z(
        \u_DataPath/pc_4_i [0]) );
  HS65_LH_AO222X4 U9929 ( .A(n7894), .B(n8689), .C(n7891), .D(
        \u_DataPath/jump_address_i [1]), .E(n8924), .F(n7889), .Z(
        \u_DataPath/pc_4_i [1]) );
  HS65_LH_AO222X4 U9930 ( .A(n7894), .B(\u_DataPath/pc_4_i [2]), .C(n7891), 
        .D(\u_DataPath/jump_address_i [2]), .E(n8923), .F(n7889), .Z(n8670) );
  HS65_LH_BFX4 U9931 ( .A(n8283), .Z(n7885) );
  HS65_LH_AO222X4 U9932 ( .A(n7894), .B(\u_DataPath/pc_4_i [3]), .C(n7891), 
        .D(\u_DataPath/jump_address_i [3]), .E(n9147), .F(n7889), .Z(n8669) );
  HS65_LH_AO222X4 U9933 ( .A(n7894), .B(\u_DataPath/pc_4_i [4]), .C(n7891), 
        .D(\u_DataPath/jump_address_i [4]), .E(n9148), .F(n7888), .Z(n8668) );
  HS65_LH_AO222X4 U9934 ( .A(n7894), .B(\u_DataPath/pc_4_i [5]), .C(n7891), 
        .D(n9409), .E(n8922), .F(n7888), .Z(n8667) );
  HS65_LH_AO222X4 U9935 ( .A(n7894), .B(\u_DataPath/pc_4_i [6]), .C(n7891), 
        .D(n9410), .E(n8921), .F(n7888), .Z(n8666) );
  HS65_LH_AO222X4 U9937 ( .A(n7894), .B(\u_DataPath/pc_4_i [7]), .C(n7891), 
        .D(\u_DataPath/jump_address_i [7]), .E(n9196), .F(n7888), .Z(n8665) );
  HS65_LH_AO222X4 U9938 ( .A(n7894), .B(\u_DataPath/pc_4_i [10]), .C(n7891), 
        .D(\u_DataPath/jump_address_i [10]), .E(n9263), .F(n7888), .Z(n8662)
         );
  HS65_LH_AO222X4 U9939 ( .A(n7894), .B(\u_DataPath/pc_4_i [8]), .C(n7891), 
        .D(n9408), .E(n8920), .F(n7888), .Z(n8664) );
  HS65_LH_AO222X4 U9940 ( .A(n7894), .B(\u_DataPath/pc_4_i [11]), .C(n7891), 
        .D(n9407), .E(n8918), .F(n7888), .Z(n8661) );
  HS65_LH_AO222X4 U9941 ( .A(n7894), .B(\u_DataPath/pc_4_i [9]), .C(n7891), 
        .D(\u_DataPath/jump_address_i [9]), .E(n9195), .F(n7888), .Z(n8663) );
  HS65_LH_AOI21X2 U9946 ( .A(n8084), .B(n8083), .C(n8117), .Z(n8085) );
  HS65_LH_CNIVX27 U9948 ( .A(rst), .Z(n8566) );
  HS65_LH_CNIVX27 U9949 ( .A(n2733), .Z(n8480) );
  HS65_LL_DFPQX4 clk_r_REG0_S1 ( .D(n2733), .CP(clk), .Q(n9334) );
  HS65_LL_DFPQX4 clk_r_REG648_S1 ( .D(Data_out_fromRAM[30]), .CP(clk), .Q(
        n9302) );
  HS65_LL_DFPQX4 clk_r_REG650_S1 ( .D(Data_out_fromRAM[29]), .CP(clk), .Q(
        n9301) );
  HS65_LL_DFPQX4 clk_r_REG652_S1 ( .D(Data_out_fromRAM[28]), .CP(clk), .Q(
        n9300) );
  HS65_LL_DFPQX4 clk_r_REG654_S1 ( .D(Data_out_fromRAM[27]), .CP(clk), .Q(
        n9299) );
  HS65_LL_DFPQX4 clk_r_REG656_S1 ( .D(Data_out_fromRAM[26]), .CP(clk), .Q(
        n9298) );
  HS65_LL_DFPQX4 clk_r_REG658_S1 ( .D(Data_out_fromRAM[25]), .CP(clk), .Q(
        n9297) );
  HS65_LL_DFPQX4 clk_r_REG663_S1 ( .D(Data_out_fromRAM[22]), .CP(clk), .Q(
        n9295) );
  HS65_LL_DFPQX4 clk_r_REG667_S1 ( .D(Data_out_fromRAM[20]), .CP(clk), .Q(
        n9293) );
  HS65_LL_DFPQX4 clk_r_REG669_S1 ( .D(Data_out_fromRAM[19]), .CP(clk), .Q(
        n9292) );
  HS65_LL_DFPQX4 clk_r_REG671_S1 ( .D(Data_out_fromRAM[18]), .CP(clk), .Q(
        n9291) );
  HS65_LL_DFPQX4 clk_r_REG673_S1 ( .D(Data_out_fromRAM[17]), .CP(clk), .Q(
        n9290) );
  HS65_LL_DFPQX4 clk_r_REG675_S1 ( .D(Data_out_fromRAM[16]), .CP(clk), .Q(
        n9289) );
  HS65_LL_DFPQX4 clk_r_REG677_S1 ( .D(Data_out_fromRAM[15]), .CP(clk), .Q(
        n9288) );
  HS65_LL_DFPQX4 clk_r_REG678_S1 ( .D(Data_out_fromRAM[14]), .CP(clk), .Q(
        n9287) );
  HS65_LL_DFPQX4 clk_r_REG679_S1 ( .D(Data_out_fromRAM[13]), .CP(clk), .Q(
        n9286) );
  HS65_LL_DFPQX4 clk_r_REG680_S1 ( .D(Data_out_fromRAM[12]), .CP(clk), .Q(
        n9285) );
  HS65_LL_DFPQX4 clk_r_REG681_S1 ( .D(Data_out_fromRAM[11]), .CP(clk), .Q(
        n9284) );
  HS65_LL_DFPQX4 clk_r_REG682_S1 ( .D(Data_out_fromRAM[10]), .CP(clk), .Q(
        n9283) );
  HS65_LL_DFPQX4 clk_r_REG683_S1 ( .D(Data_out_fromRAM[9]), .CP(clk), .Q(n9282) );
  HS65_LL_DFPQX4 clk_r_REG684_S1 ( .D(Data_out_fromRAM[8]), .CP(clk), .Q(n9281) );
  HS65_LL_DFPQX4 clk_r_REG688_S1 ( .D(Data_out_fromRAM[4]), .CP(clk), .Q(n9278) );
  HS65_LL_DFPQX4 clk_r_REG689_S1 ( .D(Data_out_fromRAM[3]), .CP(clk), .Q(n9277) );
  HS65_LL_DFPQX4 clk_r_REG690_S1 ( .D(Data_out_fromRAM[2]), .CP(clk), .Q(n9276) );
  HS65_LL_DFPQX4 clk_r_REG691_S1 ( .D(Data_out_fromRAM[1]), .CP(clk), .Q(n9275) );
  HS65_LL_DFPQX4 clk_r_REG692_S1 ( .D(Data_out_fromRAM[0]), .CP(clk), .Q(n9274) );
  HS65_LL_DFPQX4 clk_r_REG446_S2 ( .D(n7902), .CP(clk), .Q(n9272) );
  HS65_LL_DFPQX4 clk_r_REG337_S2 ( .D(\sub_x_53/A[25] ), .CP(clk), .Q(n9271)
         );
  HS65_LL_DFPQX4 clk_r_REG346_S1 ( .D(n7974), .CP(clk), .Q(n9270) );
  HS65_LL_DFPQX4 clk_r_REG389_S1 ( .D(n8001), .CP(clk), .Q(n9269) );
  HS65_LL_DFPQX4 clk_r_REG662_S1 ( .D(n8360), .CP(clk), .Q(n9268) );
  HS65_LL_DFPQX4 clk_r_REG605_S1 ( .D(n8627), .CP(clk), .Q(n9267) );
  HS65_LL_DFPQX4 clk_r_REG606_S2 ( .D(n9267), .CP(clk), .Q(n9266) );
  HS65_LL_DFPQX4 clk_r_REG173_S1 ( .D(\u_DataPath/branch_target_i [27]), .CP(
        clk), .Q(n9264) );
  HS65_LL_DFPQX4 clk_r_REG116_S1 ( .D(\u_DataPath/branch_target_i [10]), .CP(
        clk), .Q(n9263) );
  HS65_LL_DFPQX4 clk_r_REG277_S3 ( .D(n2853), .CP(clk), .Q(n9260) );
  HS65_LL_DFPQX4 clk_r_REG38_S2 ( .D(n2858), .CP(clk), .Q(n9259) );
  HS65_LL_DFPQX4 clk_r_REG406_S3 ( .D(\sub_x_53/A[30] ), .CP(clk), .Q(n9258)
         );
  HS65_LL_DFPQX4 clk_r_REG412_S2 ( .D(\sub_x_53/A[27] ), .CP(clk), .Q(n9257)
         );
  HS65_LL_DFPQX4 clk_r_REG333_S2 ( .D(\lte_x_59/B[22] ), .CP(clk), .Q(n9256)
         );
  HS65_LL_DFPQX4 clk_r_REG110_S2 ( .D(\lte_x_59/B[9] ), .CP(clk), .Q(n9255) );
  HS65_LL_DFPRQX4 clk_r_REG615_S1 ( .D(n7922), .CP(clk), .RN(n7879), .Q(n9254)
         );
  HS65_LL_DFPQX4 clk_r_REG452_S2 ( .D(n8578), .CP(clk), .Q(n9251) );
  HS65_LL_DFPQX4 clk_r_REG433_S1 ( .D(\u_DataPath/branch_target_i [0]), .CP(
        clk), .Q(n9250) );
  HS65_LL_DFPQX4 clk_r_REG374_S2 ( .D(\u_DataPath/u_execute/link_value_i [2]), 
        .CP(clk), .Q(n9249) );
  HS65_LL_DFPQX4 clk_r_REG649_S1 ( .D(n8402), .CP(clk), .Q(n9248) );
  HS65_LL_DFPQX4 clk_r_REG651_S1 ( .D(n8447), .CP(clk), .Q(n9247) );
  HS65_LL_DFPQX4 clk_r_REG661_S1 ( .D(n8370), .CP(clk), .Q(n9245) );
  HS65_LL_DFPQX4 clk_r_REG655_S1 ( .D(n8376), .CP(clk), .Q(n9244) );
  HS65_LL_DFPQX4 clk_r_REG659_S1 ( .D(n8335), .CP(clk), .Q(n9242) );
  HS65_LL_DFPQX4 clk_r_REG354_S2 ( .D(\u_DataPath/mem_writedata_out_i [28]), 
        .CP(clk), .Q(n9241) );
  HS65_LL_DFPRQX4 clk_r_REG513_S1 ( .D(n7898), .CP(clk), .RN(n9361), .Q(n9240)
         );
  HS65_LL_DFPQX4 clk_r_REG469_S4 ( .D(n7837), .CP(clk), .Q(n9239) );
  HS65_LL_DFPQX4 clk_r_REG449_S1 ( .D(\u_DataPath/cw_memwb_i [0]), .CP(clk), 
        .Q(n9238) );
  HS65_LL_DFPQX4 clk_r_REG484_S1 ( .D(\u_DataPath/cw_tomem_i [8]), .CP(clk), 
        .Q(n9237) );
  HS65_LL_DFPQX4 clk_r_REG479_S1 ( .D(\u_DataPath/cw_tomem_i [7]), .CP(clk), 
        .Q(n9236) );
  HS65_LL_DFPQX4 clk_r_REG510_S1 ( .D(\u_DataPath/cw_tomem_i [6]), .CP(clk), 
        .Q(n9235) );
  HS65_LL_DFPQX4 clk_r_REG518_S1 ( .D(\u_DataPath/cw_tomem_i [0]), .CP(clk), 
        .Q(n9234) );
  HS65_LL_DFPQX4 clk_r_REG473_S1 ( .D(\u_DataPath/jump_i ), .CP(clk), .Q(n9233) );
  HS65_LL_DFPQX4 clk_r_REG266_S1 ( .D(\u_DataPath/pc_4_to_ex_i [11]), .CP(clk), 
        .Q(n9232) );
  HS65_LL_DFPQX4 clk_r_REG259_S1 ( .D(\u_DataPath/pc_4_to_ex_i [12]), .CP(clk), 
        .Q(n9230) );
  HS65_LL_DFPQX4 clk_r_REG313_S1 ( .D(\u_DataPath/pc_4_to_ex_i [8]), .CP(clk), 
        .Q(n9229) );
  HS65_LL_DFPQX4 clk_r_REG126_S1 ( .D(\u_DataPath/pc_4_to_ex_i [13]), .CP(clk), 
        .Q(n9228) );
  HS65_LL_DFPQX4 clk_r_REG319_S1 ( .D(\u_DataPath/pc_4_to_ex_i [7]), .CP(clk), 
        .Q(n9227) );
  HS65_LL_DFPQX4 clk_r_REG132_S1 ( .D(\u_DataPath/pc_4_to_ex_i [14]), .CP(clk), 
        .Q(n9226) );
  HS65_LL_DFPQX4 clk_r_REG308_S1 ( .D(\u_DataPath/pc_4_to_ex_i [6]), .CP(clk), 
        .Q(n9225) );
  HS65_LL_DFPQX4 clk_r_REG251_S1 ( .D(\u_DataPath/pc_4_to_ex_i [15]), .CP(clk), 
        .Q(n9224) );
  HS65_LL_DFPQX4 clk_r_REG327_S1 ( .D(\u_DataPath/pc_4_to_ex_i [5]), .CP(clk), 
        .Q(n9223) );
  HS65_LL_DFPQX4 clk_r_REG244_S1 ( .D(\u_DataPath/pc_4_to_ex_i [16]), .CP(clk), 
        .Q(n9222) );
  HS65_LL_DFPQX4 clk_r_REG237_S1 ( .D(\u_DataPath/pc_4_to_ex_i [17]), .CP(clk), 
        .Q(n9221) );
  HS65_LL_DFPQX4 clk_r_REG216_S1 ( .D(\u_DataPath/pc_4_to_ex_i [18]), .CP(clk), 
        .Q(n9220) );
  HS65_LL_DFPQX4 clk_r_REG299_S1 ( .D(\u_DataPath/pc_4_to_ex_i [4]), .CP(clk), 
        .Q(n9219) );
  HS65_LL_DFPQX4 clk_r_REG224_S1 ( .D(\u_DataPath/pc_4_to_ex_i [19]), .CP(clk), 
        .Q(n9218) );
  HS65_LL_DFPQX4 clk_r_REG229_S1 ( .D(\u_DataPath/pc_4_to_ex_i [20]), .CP(clk), 
        .Q(n9217) );
  HS65_LL_DFPQX4 clk_r_REG5_S1 ( .D(\u_DataPath/pc_4_to_ex_i [3]), .CP(clk), 
        .Q(n9215) );
  HS65_LL_DFPQX4 clk_r_REG120_S1 ( .D(\u_DataPath/pc_4_to_ex_i [10]), .CP(clk), 
        .Q(n9214) );
  HS65_LL_DFPQX4 clk_r_REG156_S1 ( .D(\u_DataPath/pc_4_to_ex_i [22]), .CP(clk), 
        .Q(n9213) );
  HS65_LL_DFPQX4 clk_r_REG367_S1 ( .D(\u_DataPath/u_execute/link_value_i [1]), 
        .CP(clk), .Q(n9212) );
  HS65_LL_DFPQX4 clk_r_REG209_S1 ( .D(\u_DataPath/pc_4_to_ex_i [23]), .CP(clk), 
        .Q(n9210) );
  HS65_LL_DFPQX4 clk_r_REG161_S1 ( .D(\u_DataPath/pc_4_to_ex_i [24]), .CP(clk), 
        .Q(n9209) );
  HS65_LL_DFPQX4 clk_r_REG166_S1 ( .D(\u_DataPath/pc_4_to_ex_i [25]), .CP(clk), 
        .Q(n9208) );
  HS65_LL_DFPQX4 clk_r_REG171_S1 ( .D(\u_DataPath/pc_4_to_ex_i [26]), .CP(clk), 
        .Q(n9207) );
  HS65_LL_DFPQX4 clk_r_REG177_S1 ( .D(\u_DataPath/pc_4_to_ex_i [27]), .CP(clk), 
        .Q(n9206) );
  HS65_LL_DFPQX4 clk_r_REG183_S1 ( .D(\u_DataPath/pc_4_to_ex_i [28]), .CP(clk), 
        .Q(n9205) );
  HS65_LL_DFPQX4 clk_r_REG200_S1 ( .D(\u_DataPath/pc_4_to_ex_i [29]), .CP(clk), 
        .Q(n9204) );
  HS65_LL_DFPQX4 clk_r_REG188_S1 ( .D(\u_DataPath/pc_4_to_ex_i [30]), .CP(clk), 
        .Q(n9203) );
  HS65_LL_DFPQX4 clk_r_REG193_S1 ( .D(\u_DataPath/pc_4_to_ex_i [31]), .CP(clk), 
        .Q(n9202) );
  HS65_LL_DFPQX4 clk_r_REG343_S3 ( .D(\lte_x_59/B[15] ), .CP(clk), .Q(n9200)
         );
  HS65_LL_DFPQX4 clk_r_REG203_S1 ( .D(\u_DataPath/branch_target_i [25]), .CP(
        clk), .Q(n9199) );
  HS65_LL_DFPQX4 clk_r_REG128_S1 ( .D(\u_DataPath/branch_target_i [14]), .CP(
        clk), .Q(n9198) );
  HS65_LL_DFPQX4 clk_r_REG210_S1 ( .D(\u_DataPath/branch_target_i [23]), .CP(
        clk), .Q(n9197) );
  HS65_LL_DFPQX4 clk_r_REG315_S1 ( .D(\u_DataPath/branch_target_i [7]), .CP(
        clk), .Q(n9196) );
  HS65_LL_DFPQX4 clk_r_REG240_S1 ( .D(\u_DataPath/branch_target_i [16]), .CP(
        clk), .Q(n9194) );
  HS65_LL_DFPQX4 clk_r_REG135_S1 ( .D(\u_DataPath/branch_target_i [21]), .CP(
        clk), .Q(n9193) );
  HS65_LL_DFPRQX4 clk_r_REG535_S1 ( .D(n7921), .CP(clk), .RN(n9354), .Q(n9191)
         );
  HS65_LL_DFPQX4 clk_r_REG468_S4 ( .D(n7904), .CP(clk), .Q(n9190) );
  HS65_LL_DFPQX4 clk_r_REG471_S4 ( .D(n7903), .CP(clk), .Q(n9189) );
  HS65_LL_DFPQX4 clk_r_REG462_S1 ( .D(n7882), .CP(clk), .Q(n9188) );
  HS65_LL_DFPQX4 clk_r_REG472_S4 ( .D(n7907), .CP(clk), .Q(n9187) );
  HS65_LL_DFPQX4 clk_r_REG602_S1 ( .D(n8629), .CP(clk), .Q(n9185) );
  HS65_LL_DFPQX4 clk_r_REG603_S2 ( .D(n9185), .CP(clk), .Q(n9184) );
  HS65_LL_DFPQX4 clk_r_REG599_S1 ( .D(n8631), .CP(clk), .Q(n9183) );
  HS65_LL_DFPQX4 clk_r_REG600_S2 ( .D(n9183), .CP(clk), .Q(n9182) );
  HS65_LL_DFPQX4 clk_r_REG608_S1 ( .D(n8623), .CP(clk), .Q(n9181) );
  HS65_LL_DFPQX4 clk_r_REG609_S2 ( .D(n9181), .CP(clk), .Q(n9180) );
  HS65_LL_DFPQX4 clk_r_REG588_S1 ( .D(\u_DataPath/u_idexreg/N31 ), .CP(clk), 
        .Q(n9179) );
  HS65_LL_DFPQX4 clk_r_REG545_S1 ( .D(\u_DataPath/u_idexreg/N33 ), .CP(clk), 
        .Q(n9177) );
  HS65_LL_DFPQX4 clk_r_REG546_S2 ( .D(n9177), .CP(clk), .Q(n9176) );
  HS65_LL_DFPQX4 clk_r_REG542_S1 ( .D(\u_DataPath/immediate_ext_ex_i [7]), 
        .CP(clk), .Q(n9175) );
  HS65_LL_DFPQX4 clk_r_REG543_S2 ( .D(n9175), .CP(clk), .Q(n9174) );
  HS65_LL_DFPQX4 clk_r_REG548_S1 ( .D(\u_DataPath/immediate_ext_ex_i [9]), 
        .CP(clk), .Q(n9173) );
  HS65_LL_DFPQX4 clk_r_REG549_S2 ( .D(n9173), .CP(clk), .Q(n9172) );
  HS65_LL_DFPQX4 clk_r_REG552_S2 ( .D(n9171), .CP(clk), .Q(n9170) );
  HS65_LL_DFPQX4 clk_r_REG571_S3 ( .D(n8162), .CP(clk), .Q(n9169) );
  HS65_LL_DFPQX4 clk_r_REG527_S2 ( .D(n8070), .CP(clk), .Q(n9168) );
  HS65_LL_DFPQX4 clk_r_REG509_S3 ( .D(n8055), .CP(clk), .Q(n9167) );
  HS65_LL_DFPQX4 clk_r_REG685_S1 ( .D(n8302), .CP(clk), .Q(n9166) );
  HS65_LL_DFPQX4 clk_r_REG194_S1 ( .D(\u_DataPath/branch_target_i [31]), .CP(
        clk), .Q(n9165) );
  HS65_LL_DFPQX4 clk_r_REG201_S1 ( .D(\u_DataPath/branch_target_i [29]), .CP(
        clk), .Q(n9164) );
  HS65_LL_DFPRQX4 clk_r_REG555_S2 ( .D(n7918), .CP(clk), .RN(n9356), .Q(n9153)
         );
  HS65_LL_DFPQX4 clk_r_REG442_S3 ( .D(n8054), .CP(clk), .Q(n9152) );
  HS65_LL_DFPQX4 clk_r_REG464_S3 ( .D(\u_DataPath/cw_exmem_i [9]), .CP(clk), 
        .Q(n9151) );
  HS65_LL_DFPQX4 clk_r_REG385_S3 ( .D(n8271), .CP(clk), .Q(n9150) );
  HS65_LL_DFPQX4 clk_r_REG489_S3 ( .D(n8095), .CP(clk), .Q(n9149) );
  HS65_LL_DFPQX4 clk_r_REG322_S1 ( .D(\u_DataPath/branch_target_i [4]), .CP(
        clk), .Q(n9148) );
  HS65_LL_DFPQX4 clk_r_REG611_S1 ( .D(n8625), .CP(clk), .Q(n9145) );
  HS65_LL_DFPQX4 clk_r_REG612_S2 ( .D(n9145), .CP(clk), .Q(n9144) );
  HS65_LL_DFPRQX4 clk_r_REG538_S2 ( .D(n7920), .CP(clk), .RN(n9355), .Q(n9141)
         );
  HS65_LL_DFPQX4 clk_r_REG448_S2 ( .D(n7914), .CP(clk), .Q(n9140) );
  HS65_LL_DFPRQX4 clk_r_REG514_S1 ( .D(n7924), .CP(clk), .RN(n9354), .Q(n9138)
         );
  HS65_LL_DFPQX4 clk_r_REG470_S4 ( .D(n7849), .CP(clk), .Q(n9137) );
  HS65_LL_DFPQX4 clk_r_REG461_S1 ( .D(n7881), .CP(clk), .Q(n9136) );
  HS65_LL_DFPQX4 clk_r_REG467_S1 ( .D(n7908), .CP(clk), .Q(n9135) );
  HS65_LL_DFPQX4 clk_r_REG460_S1 ( .D(n7883), .CP(clk), .Q(n9134) );
  HS65_LL_DFPQX4 clk_r_REG459_S1 ( .D(n7884), .CP(clk), .Q(n9133) );
  HS65_LL_DFPRQX4 clk_r_REG511_S1 ( .D(n7897), .CP(clk), .RN(n9355), .Q(n9131)
         );
  HS65_LL_DFPQX4 clk_r_REG647_S1 ( .D(n8420), .CP(clk), .Q(n9129) );
  HS65_LL_DFPQX4 clk_r_REG383_S3 ( .D(n8299), .CP(clk), .Q(n9127) );
  HS65_LL_DFPQX4 clk_r_REG666_S1 ( .D(n8365), .CP(clk), .Q(n9126) );
  HS65_LL_DFPQX4 clk_r_REG672_S1 ( .D(n8454), .CP(clk), .Q(n9125) );
  HS65_LL_DFPQX4 clk_r_REG670_S1 ( .D(n8324), .CP(clk), .Q(n9124) );
  HS65_LL_DFPQX4 clk_r_REG664_S1 ( .D(n8351), .CP(clk), .Q(n9123) );
  HS65_LL_DFPQX4 clk_r_REG676_S1 ( .D(n8356), .CP(clk), .Q(n9122) );
  HS65_LL_DFPQX4 clk_r_REG674_S1 ( .D(n8406), .CP(clk), .Q(n9121) );
  HS65_LL_DFPQX4 clk_r_REG668_S1 ( .D(n8410), .CP(clk), .Q(n9120) );
  HS65_LL_DFPQX4 clk_r_REG447_S1 ( .D(n7899), .CP(clk), .Q(n9119) );
  HS65_LL_DFPQX4 clk_r_REG45_S1 ( .D(\u_DataPath/u_execute/psw_status_i [1]), 
        .CP(clk), .Q(n9118) );
  HS65_LL_DFPQX4 clk_r_REG373_S1 ( .D(\u_DataPath/pc_4_to_ex_i [2]), .CP(clk), 
        .Q(n9116) );
  HS65_LL_DFPQX4 clk_r_REG430_S1 ( .D(\u_DataPath/u_execute/link_value_i [0]), 
        .CP(clk), .Q(n9115) );
  HS65_LL_DFPQX4 clk_r_REG444_S1 ( .D(\u_DataPath/reg_write_i ), .CP(clk), .Q(
        n9111) );
  HS65_LL_DFPQX4 clk_r_REG465_S1 ( .D(\u_DataPath/cw_memwb_i [1]), .CP(clk), 
        .Q(n9110) );
  HS65_LL_DFPQX4 clk_r_REG458_S1 ( .D(n7885), .CP(clk), .Q(n9109) );
  HS65_LL_DFPRQX4 clk_r_REG191_S4 ( .D(\u_DataPath/pc_4_i [31]), .CP(clk), 
        .RN(n9361), .Q(n9108) );
  HS65_LL_DFPQX4 clk_r_REG68_S2 ( .D(\sub_x_53/A[29] ), .CP(clk), .Q(n9107) );
  HS65_LL_DFPQX4 clk_r_REG26_S3 ( .D(\lte_x_59/B[18] ), .CP(clk), .Q(n9106) );
  HS65_LL_DFPQX4 clk_r_REG52_S2 ( .D(\lte_x_59/B[1] ), .CP(clk), .Q(n9105) );
  HS65_LL_DFPQX4 clk_r_REG350_S2 ( .D(n3474), .CP(clk), .Q(n9104) );
  HS65_LL_DFPQX4 clk_r_REG394_S3 ( .D(n8575), .CP(clk), .Q(n9103) );
  HS65_LL_DFPQX4 clk_r_REG594_S3 ( .D(n8076), .CP(clk), .Q(n9102) );
  HS65_LL_DFPQX4 clk_r_REG134_S2 ( .D(\u_DataPath/u_execute/link_value_i [14]), 
        .CP(clk), .Q(n9101) );
  HS65_LL_DFPQX4 clk_r_REG301_S2 ( .D(\u_DataPath/u_execute/link_value_i [7]), 
        .CP(clk), .Q(n9100) );
  HS65_LL_DFPQX4 clk_r_REG581_S3 ( .D(n8115), .CP(clk), .Q(n9099) );
  HS65_LL_DFPQX4 clk_r_REG347_S3 ( .D(n2842), .CP(clk), .Q(n9096) );
  HS65_LL_DFPQX4 clk_r_REG92_S2 ( .D(\sub_x_53/A[17] ), .CP(clk), .Q(n9094) );
  HS65_LL_DFPQX4 clk_r_REG417_S2 ( .D(\lte_x_59/B[16] ), .CP(clk), .Q(n9093)
         );
  HS65_LL_DFPQX4 clk_r_REG10_S3 ( .D(\sub_x_53/A[0] ), .CP(clk), .Q(n9092) );
  HS65_LL_DFPQX4 clk_r_REG403_S4 ( .D(\lte_x_59/B[8] ), .CP(clk), .Q(n9091) );
  HS65_LL_DFPQX4 clk_r_REG32_S3 ( .D(n7867), .CP(clk), .Q(n9090) );
  HS65_LL_DFPQX4 clk_r_REG107_S4 ( .D(\lte_x_59/B[21] ), .CP(clk), .Q(n9089)
         );
  HS65_LL_DFPQX4 clk_r_REG421_S3 ( .D(n3521), .CP(clk), .Q(n9088) );
  HS65_LL_DFPRQX4 clk_r_REG181_S4 ( .D(\u_DataPath/pc_4_i [28]), .CP(clk), 
        .RN(n8677), .Q(n9087) );
  HS65_LL_DFPQX4 clk_r_REG384_S3 ( .D(n8452), .CP(clk), .Q(n9086) );
  HS65_LL_DFPQX4 clk_r_REG339_S1 ( .D(\u_DataPath/mem_writedata_out_i [25]), 
        .CP(clk), .Q(n9085) );
  HS65_LL_DFPQX4 clk_r_REG508_S3 ( .D(n9084), .CP(clk), .Q(n9083) );
  HS65_LL_DFPQX4 clk_r_REG375_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [3]), 
        .CP(clk), .Q(n9080) );
  HS65_LL_DFPQX4 clk_r_REG303_S2 ( .D(\u_DataPath/u_execute/link_value_i [6]), 
        .CP(clk), .Q(n9079) );
  HS65_LL_DFPQX4 clk_r_REG503_S1 ( .D(\u_DataPath/regfile_addr_out_towb_i [2]), 
        .CP(clk), .Q(n9078) );
  HS65_LL_DFPQX4 clk_r_REG530_S1 ( .D(\u_DataPath/idex_rt_i [3]), .CP(clk), 
        .Q(n9077) );
  HS65_LL_DFPQX4 clk_r_REG501_S1 ( .D(\u_DataPath/regfile_addr_out_towb_i [0]), 
        .CP(clk), .Q(n9076) );
  HS65_LL_DFPQX4 clk_r_REG497_S1 ( .D(\u_DataPath/regfile_addr_out_towb_i [3]), 
        .CP(clk), .Q(n9075) );
  HS65_LL_DFPQX4 clk_r_REG85_S2 ( .D(n7855), .CP(clk), .Q(n9074) );
  HS65_LL_DFPQX4 clk_r_REG79_S3 ( .D(n8458), .CP(clk), .Q(n9073) );
  HS65_LL_DFPQX4 clk_r_REG108_S2 ( .D(n8474), .CP(clk), .Q(n9072) );
  HS65_LL_DFPQX4 clk_r_REG100_S3 ( .D(\sub_x_53/A[23] ), .CP(clk), .Q(n9071)
         );
  HS65_LL_DFPRQX4 clk_r_REG175_S3 ( .D(\u_DataPath/pc_4_i [27]), .CP(clk), 
        .RN(n9361), .Q(n9070) );
  HS65_LL_DFPQX4 clk_r_REG246_S2 ( .D(n7865), .CP(clk), .Q(n9065) );
  HS65_LL_DFPQX4 clk_r_REG93_S2 ( .D(n7857), .CP(clk), .Q(n9063) );
  HS65_LL_DFPQX4 clk_r_REG24_S2 ( .D(n7842), .CP(clk), .Q(n9062) );
  HS65_LL_DFPQX4 clk_r_REG20_S2 ( .D(n7850), .CP(clk), .Q(n9061) );
  HS65_LL_DFPQX4 clk_r_REG104_S3 ( .D(n7844), .CP(clk), .Q(n9060) );
  HS65_LL_DFPQX4 clk_r_REG95_S3 ( .D(n8471), .CP(clk), .Q(n9059) );
  HS65_LL_DFPQX4 clk_r_REG87_S2 ( .D(n8466), .CP(clk), .Q(n9058) );
  HS65_LL_DFPQX4 clk_r_REG97_S4 ( .D(\sub_x_53/A[20] ), .CP(clk), .Q(n9056) );
  HS65_LL_DFPQX4 clk_r_REG340_S4 ( .D(\lte_x_59/B[24] ), .CP(clk), .Q(n9055)
         );
  HS65_LL_DFPQX4 clk_r_REG167_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [26]), 
        .CP(clk), .Q(n9054) );
  HS65_LL_DFPQX4 clk_r_REG8_S2 ( .D(\lte_x_59/B[3] ), .CP(clk), .Q(n9053) );
  HS65_LL_DFPQX4 clk_r_REG517_S2 ( .D(n8636), .CP(clk), .Q(n9052) );
  HS65_LL_DFPQX4 clk_r_REG393_S3 ( .D(n8300), .CP(clk), .Q(n9051) );
  HS65_LL_DFPQX4 clk_r_REG483_S3 ( .D(n8068), .CP(clk), .Q(n9050) );
  HS65_LL_DFPQX4 clk_r_REG477_S3 ( .D(n8069), .CP(clk), .Q(n9049) );
  HS65_LL_DFPQX4 clk_r_REG456_S3 ( .D(n8634), .CP(clk), .Q(n9048) );
  HS65_LL_DFPQX4 clk_r_REG218_S2 ( .D(n5703), .CP(clk), .Q(n9047) );
  HS65_LL_DFPQX4 clk_r_REG219_S2 ( .D(\u_DataPath/u_execute/link_value_i [20]), 
        .CP(clk), .Q(n9046) );
  HS65_LL_DFPQX4 clk_r_REG115_S2 ( .D(\u_DataPath/u_execute/link_value_i [9]), 
        .CP(clk), .Q(n9045) );
  HS65_LL_DFPQX4 clk_r_REG260_S2 ( .D(\u_DataPath/u_execute/link_value_i [12]), 
        .CP(clk), .Q(n9044) );
  HS65_LL_DFPQX4 clk_r_REG267_S2 ( .D(n4006), .CP(clk), .Q(n9043) );
  HS65_LL_DFPQX4 clk_r_REG330_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [4]), 
        .CP(clk), .Q(n9041) );
  HS65_LL_DFPQX4 clk_r_REG328_S2 ( .D(\u_DataPath/u_execute/link_value_i [5]), 
        .CP(clk), .Q(n9040) );
  HS65_LL_DFPQX4 clk_r_REG567_S1 ( .D(\u_DataPath/immediate_ext_ex_i [2]), 
        .CP(clk), .Q(n9039) );
  HS65_LL_DFPQX4 clk_r_REG568_S2 ( .D(n9039), .CP(clk), .Q(n9038) );
  HS65_LL_DFPQX4 clk_r_REG579_S1 ( .D(\u_DataPath/immediate_ext_ex_i [1]), 
        .CP(clk), .Q(n9037) );
  HS65_LL_DFPQX4 clk_r_REG580_S2 ( .D(n9037), .CP(clk), .Q(n9036) );
  HS65_LL_DFPQX4 clk_r_REG586_S2 ( .D(n9035), .CP(clk), .Q(n9034) );
  HS65_LL_DFPQX4 clk_r_REG574_S1 ( .D(\u_DataPath/immediate_ext_ex_i [3]), 
        .CP(clk), .Q(n9033) );
  HS65_LL_DFPQX4 clk_r_REG575_S2 ( .D(n9033), .CP(clk), .Q(n9032) );
  HS65_LL_DFPQX4 clk_r_REG505_S1 ( .D(\u_DataPath/regfile_addr_out_towb_i [1]), 
        .CP(clk), .Q(n9031) );
  HS65_LL_DFPQX4 clk_r_REG592_S1 ( .D(\u_DataPath/immediate_ext_ex_i [5]), 
        .CP(clk), .Q(n9030) );
  HS65_LL_DFPQX4 clk_r_REG593_S2 ( .D(n9030), .CP(clk), .Q(n9029) );
  HS65_LL_DFPQX4 clk_r_REG73_S2 ( .D(n8477), .CP(clk), .Q(n9028) );
  HS65_LL_DFPQX4 clk_r_REG63_S2 ( .D(n8469), .CP(clk), .Q(n9026) );
  HS65_LL_DFPQX4 clk_r_REG195_S1 ( .D(\u_DataPath/branch_target_i [30]), .CP(
        clk), .Q(n9025) );
  HS65_LL_DFPQX4 clk_r_REG196_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [29]), 
        .CP(clk), .Q(n9024) );
  HS65_LL_DFPQX4 clk_r_REG178_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [27]), 
        .CP(clk), .Q(n9023) );
  HS65_LL_DFPQX4 clk_r_REG19_S2 ( .D(\lte_x_59/B[14] ), .CP(clk), .Q(n9022) );
  HS65_LL_DFPQX4 clk_r_REG41_S3 ( .D(\sub_x_53/A[2] ), .CP(clk), .Q(n9021) );
  HS65_LL_DFPQX4 clk_r_REG34_S1 ( .D(\u_DataPath/mem_writedata_out_i [8]), 
        .CP(clk), .Q(n9019) );
  HS65_LL_DFPQX4 clk_r_REG388_S3 ( .D(\u_DataPath/mem_writedata_out_i [0]), 
        .CP(clk), .Q(n9018) );
  HS65_LL_DFPQX4 clk_r_REG238_S2 ( .D(\u_DataPath/u_execute/link_value_i [17]), 
        .CP(clk), .Q(n9017) );
  HS65_LL_DFPQX4 clk_r_REG463_S3 ( .D(n8059), .CP(clk), .Q(n9016) );
  HS65_LL_DFPQX4 clk_r_REG127_S2 ( .D(\u_DataPath/u_execute/link_value_i [13]), 
        .CP(clk), .Q(n9015) );
  HS65_LL_DFPQX4 clk_r_REG133_S2 ( .D(\u_DataPath/u_execute/link_value_i [15]), 
        .CP(clk), .Q(n9014) );
  HS65_LL_DFPQX4 clk_r_REG271_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [9]), 
        .CP(clk), .Q(n9013) );
  HS65_LL_DFPQX4 clk_r_REG616_S1 ( .D(n8117), .CP(clk), .Q(n9012) );
  HS65_LL_DFPQX4 clk_r_REG320_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [7]), 
        .CP(clk), .Q(n9011) );
  HS65_LL_DFPQX4 clk_r_REG300_S2 ( .D(\u_DataPath/u_execute/link_value_i [4]), 
        .CP(clk), .Q(n9008) );
  HS65_LL_DFPQX4 clk_r_REG6_S2 ( .D(\u_DataPath/u_execute/link_value_i [3]), 
        .CP(clk), .Q(n9006) );
  HS65_LL_DFPQX4 clk_r_REG566_S3 ( .D(n8121), .CP(clk), .Q(n9005) );
  HS65_LL_DFPQX4 clk_r_REG558_S1 ( .D(\u_DataPath/rs_ex_i [3]), .CP(clk), .Q(
        n9004) );
  HS65_LL_DFPQX4 clk_r_REG572_S3 ( .D(n8096), .CP(clk), .Q(n9003) );
  HS65_LL_DFPQX4 clk_r_REG30_S2 ( .D(n7859), .CP(clk), .Q(n9001) );
  HS65_LL_DFPQX4 clk_r_REG148_S2 ( .D(\u_DataPath/u_execute/link_value_i [31]), 
        .CP(clk), .Q(n9000) );
  HS65_LL_DFPQX4 clk_r_REG184_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [30]), 
        .CP(clk), .Q(n8999) );
  HS65_LL_DFPQX4 clk_r_REG179_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [28]), 
        .CP(clk), .Q(n8998) );
  HS65_LL_DFPQX4 clk_r_REG425_S2 ( .D(\lte_x_59/B[7] ), .CP(clk), .Q(n8997) );
  HS65_LL_DFPQX4 clk_r_REG145_S2 ( .D(\u_DataPath/u_execute/link_value_i [27]), 
        .CP(clk), .Q(n8996) );
  HS65_LL_DFPRQX4 clk_r_REG159_S4 ( .D(\u_DataPath/pc_4_i [24]), .CP(clk), 
        .RN(n8677), .Q(n8992) );
  HS65_LL_DFPRQX4 clk_r_REG137_S3 ( .D(\u_DataPath/pc_4_i [21]), .CP(clk), 
        .RN(n9354), .Q(n8991) );
  HS65_LL_DFPQX4 clk_r_REG162_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [25]), 
        .CP(clk), .Q(n8990) );
  HS65_LL_DFPRQX4 clk_r_REG207_S4 ( .D(\u_DataPath/pc_4_i [23]), .CP(clk), 
        .RN(n9361), .Q(n8989) );
  HS65_LL_DFPQX4 clk_r_REG144_S2 ( .D(\u_DataPath/u_execute/link_value_i [25]), 
        .CP(clk), .Q(n8987) );
  HS65_LL_DFPRQX4 clk_r_REG242_S3 ( .D(\u_DataPath/pc_4_i [16]), .CP(clk), 
        .RN(n8677), .Q(n8986) );
  HS65_LL_DFPRQX4 clk_r_REG227_S3 ( .D(\u_DataPath/pc_4_i [20]), .CP(clk), 
        .RN(n9361), .Q(n8985) );
  HS65_LL_DFPQX4 clk_r_REG143_S2 ( .D(\u_DataPath/u_execute/link_value_i [24]), 
        .CP(clk), .Q(n8983) );
  HS65_LL_DFPQX4 clk_r_REG231_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [19]), 
        .CP(clk), .Q(n8982) );
  HS65_LL_DFPRQX4 clk_r_REG124_S3 ( .D(\u_DataPath/pc_4_i [13]), .CP(clk), 
        .RN(n9361), .Q(n8981) );
  HS65_LL_DFPRQX4 clk_r_REG264_S3 ( .D(\u_DataPath/pc_4_i [11]), .CP(clk), 
        .RN(n9361), .Q(n8978) );
  HS65_LL_DFPQX4 clk_r_REG205_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [23]), 
        .CP(clk), .Q(n8977) );
  HS65_LL_DFPQX4 clk_r_REG142_S2 ( .D(\u_DataPath/u_execute/link_value_i [23]), 
        .CP(clk), .Q(n8975) );
  HS65_LL_DFPRQX4 clk_r_REG118_S3 ( .D(\u_DataPath/pc_4_i [10]), .CP(clk), 
        .RN(n2877), .Q(n8974) );
  HS65_LL_DFPQX4 clk_r_REG217_S2 ( .D(n4288), .CP(clk), .Q(n8972) );
  HS65_LL_DFPQX4 clk_r_REG522_S1 ( .D(\u_DataPath/rs_ex_i [0]), .CP(clk), .Q(
        n8969) );
  HS65_LL_DFPQX4 clk_r_REG524_S1 ( .D(\u_DataPath/idex_rt_i [4]), .CP(clk), 
        .Q(n8968) );
  HS65_LL_DFPQX4 clk_r_REG554_S1 ( .D(\u_DataPath/idex_rt_i [2]), .CP(clk), 
        .Q(n8967) );
  HS65_LL_DFPQX4 clk_r_REG532_S1 ( .D(\u_DataPath/idex_rt_i [1]), .CP(clk), 
        .Q(n8966) );
  HS65_LL_DFPQX4 clk_r_REG578_S3 ( .D(n8092), .CP(clk), .Q(n8965) );
  HS65_LL_DFPQX4 clk_r_REG565_S3 ( .D(n8089), .CP(clk), .Q(n8964) );
  HS65_LL_DFPRQX4 clk_r_REG306_S3 ( .D(\u_DataPath/pc_4_i [6]), .CP(clk), .RN(
        n9361), .Q(n8963) );
  HS65_LL_DFPRQX4 clk_r_REG214_S3 ( .D(\u_DataPath/pc_4_i [18]), .CP(clk), 
        .RN(n2877), .Q(n8962) );
  HS65_LL_DFPQX4 clk_r_REG443_S1 ( .D(n7833), .CP(clk), .Q(n8961) );
  HS65_LL_DFPQX4 clk_r_REG499_S1 ( .D(\u_DataPath/regfile_addr_out_towb_i [4]), 
        .CP(clk), .Q(n8960) );
  HS65_LL_DFPQX4 clk_r_REG232_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [18]), 
        .CP(clk), .Q(n8958) );
  HS65_LL_DFPQX4 clk_r_REG239_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [17]), 
        .CP(clk), .Q(n8957) );
  HS65_LL_DFPQX4 clk_r_REG230_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [20]), 
        .CP(clk), .Q(n8956) );
  HS65_LL_DFPQX4 clk_r_REG314_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [8]), 
        .CP(clk), .Q(n8955) );
  HS65_LL_DFPQX4 clk_r_REG329_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [5]), 
        .CP(clk), .Q(n8954) );
  HS65_LL_DFPQX4 clk_r_REG151_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [21]), 
        .CP(clk), .Q(n8953) );
  HS65_LL_DFPQX4 clk_r_REG254_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [13]), 
        .CP(clk), .Q(n8952) );
  HS65_LL_DFPQX4 clk_r_REG269_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [10]), 
        .CP(clk), .Q(n8951) );
  HS65_LL_DFPQX4 clk_r_REG252_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [15]), 
        .CP(clk), .Q(n8949) );
  HS65_LL_DFPQX4 clk_r_REG253_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [14]), 
        .CP(clk), .Q(n8948) );
  HS65_LL_DFPQX4 clk_r_REG302_S2 ( .D(\u_DataPath/u_execute/link_value_i [8]), 
        .CP(clk), .Q(n8947) );
  HS65_LL_DFPQX4 clk_r_REG245_S2 ( .D(n5690), .CP(clk), .Q(n8946) );
  HS65_LL_DFPQX4 clk_r_REG369_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [2]), 
        .CP(clk), .Q(n8945) );
  HS65_LL_DFPQX4 clk_r_REG560_S1 ( .D(\u_DataPath/rs_ex_i [1]), .CP(clk), .Q(
        n8944) );
  HS65_LL_DFPQX4 clk_r_REG520_S1 ( .D(\u_DataPath/rs_ex_i [2]), .CP(clk), .Q(
        n8943) );
  HS65_LL_DFPQX4 clk_r_REG534_S1 ( .D(\u_DataPath/idex_rt_i [0]), .CP(clk), 
        .Q(n8942) );
  HS65_LL_DFPQX4 clk_r_REG202_S1 ( .D(\u_DataPath/branch_target_i [28]), .CP(
        clk), .Q(n8941) );
  HS65_LL_DFPQX4 clk_r_REG172_S1 ( .D(\u_DataPath/branch_target_i [26]), .CP(
        clk), .Q(n8940) );
  HS65_LL_DFPQX4 clk_r_REG140_S2 ( .D(n5169), .CP(clk), .Q(n8939) );
  HS65_LL_DFPQX4 clk_r_REG141_S2 ( .D(n5698), .CP(clk), .Q(n8938) );
  HS65_LL_DFPQX4 clk_r_REG432_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [0]), 
        .CP(clk), .Q(n8937) );
  HS65_LL_DFPQX4 clk_r_REG189_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [31]), 
        .CP(clk), .Q(n8936) );
  HS65_LL_DFPQX4 clk_r_REG157_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [24]), 
        .CP(clk), .Q(n8934) );
  HS65_LL_DFPQX4 clk_r_REG152_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [22]), 
        .CP(clk), .Q(n8933) );
  HS65_LL_DFPQX4 clk_r_REG453_S1 ( .D(
        \u_DataPath/u_decode_unit/hdu_0/current_state [1]), .CP(clk), .Q(n8932) );
  HS65_LL_DFPQX4 clk_r_REG204_S1 ( .D(\u_DataPath/branch_target_i [24]), .CP(
        clk), .Q(n8931) );
  HS65_LL_DFPQX4 clk_r_REG247_S1 ( .D(\u_DataPath/branch_target_i [15]), .CP(
        clk), .Q(n8930) );
  HS65_LL_DFPQX4 clk_r_REG233_S1 ( .D(\u_DataPath/branch_target_i [17]), .CP(
        clk), .Q(n8928) );
  HS65_LL_DFPQX4 clk_r_REG212_S1 ( .D(\u_DataPath/branch_target_i [18]), .CP(
        clk), .Q(n8927) );
  HS65_LL_DFPQX4 clk_r_REG225_S1 ( .D(\u_DataPath/branch_target_i [20]), .CP(
        clk), .Q(n8926) );
  HS65_LL_DFPQX4 clk_r_REG220_S1 ( .D(\u_DataPath/branch_target_i [19]), .CP(
        clk), .Q(n8925) );
  HS65_LL_DFPQX4 clk_r_REG379_S1 ( .D(\u_DataPath/branch_target_i [1]), .CP(
        clk), .Q(n8924) );
  HS65_LL_DFPQX4 clk_r_REG376_S1 ( .D(\u_DataPath/branch_target_i [2]), .CP(
        clk), .Q(n8923) );
  HS65_LL_DFPQX4 clk_r_REG323_S1 ( .D(\u_DataPath/branch_target_i [5]), .CP(
        clk), .Q(n8922) );
  HS65_LL_DFPQX4 clk_r_REG304_S1 ( .D(\u_DataPath/branch_target_i [6]), .CP(
        clk), .Q(n8921) );
  HS65_LL_DFPQX4 clk_r_REG309_S1 ( .D(\u_DataPath/branch_target_i [8]), .CP(
        clk), .Q(n8920) );
  HS65_LL_DFPQX4 clk_r_REG262_S1 ( .D(\u_DataPath/branch_target_i [11]), .CP(
        clk), .Q(n8918) );
  HS65_LL_DFPQX4 clk_r_REG255_S1 ( .D(\u_DataPath/branch_target_i [12]), .CP(
        clk), .Q(n8917) );
  HS65_LL_DFPQX4 clk_r_REG441_S3 ( .D(n8053), .CP(clk), .Q(n8916) );
  HS65_LL_DFPQX4 clk_r_REG62_S1 ( .D(\u_DataPath/from_alu_data_out_i [28]), 
        .CP(clk), .Q(n8914) );
  HS65_LL_DFPQX4 clk_r_REG596_S1 ( .D(\u_DataPath/immediate_ext_ex_i [4]), 
        .CP(clk), .Q(n8913) );
  HS65_LL_DFPQX4 clk_r_REG597_S2 ( .D(n8913), .CP(clk), .Q(n8912) );
  HS65_LL_DFPQX4 clk_r_REG457_S3 ( .D(\u_DataPath/cw_to_ex_i [20]), .CP(clk), 
        .Q(n8910) );
  HS65_LL_DFPQX4 clk_r_REG77_S1 ( .D(\u_DataPath/from_alu_data_out_i [15]), 
        .CP(clk), .Q(n8909) );
  HS65_LL_DFPQX4 clk_r_REG71_S1 ( .D(\u_DataPath/from_alu_data_out_i [10]), 
        .CP(clk), .Q(n8907) );
  HS65_LL_DFPQX4 clk_r_REG445_S2 ( .D(n7306), .CP(clk), .Q(n8906) );
  HS65_LL_DFPQX4 clk_r_REG355_S2 ( .D(\lte_x_59/B[28] ), .CP(clk), .Q(n8905)
         );
  HS65_LL_DFPQX4 clk_r_REG47_S3 ( .D(\u_DataPath/dataOut_exe_i [1]), .CP(clk), 
        .Q(n8904) );
  HS65_LL_DFPQX4 clk_r_REG58_S4 ( .D(n8465), .CP(clk), .Q(n8903) );
  HS65_LL_DFPQX4 clk_r_REG27_S3 ( .D(n8461), .CP(clk), .Q(n8902) );
  HS65_LL_DFPQX4 clk_r_REG82_S2 ( .D(n8478), .CP(clk), .Q(n8900) );
  HS65_LL_DFPQX4 clk_r_REG42_S3 ( .D(n7841), .CP(clk), .Q(n8899) );
  HS65_LL_DFPQX4 clk_r_REG391_S3 ( .D(n8301), .CP(clk), .Q(n8898) );
  HS65_LL_DFPQX4 clk_r_REG392_S3 ( .D(n8318), .CP(clk), .Q(n8897) );
  HS65_LL_DFPQX4 clk_r_REG9_S2 ( .D(n7860), .CP(clk), .Q(n8896) );
  HS65_LL_DFPQX4 clk_r_REG17_S2 ( .D(n8475), .CP(clk), .Q(n8895) );
  HS65_LL_DFPQX4 clk_r_REG53_S3 ( .D(n8463), .CP(clk), .Q(n8893) );
  HS65_LL_DFPQX4 clk_r_REG476_S3 ( .D(n8128), .CP(clk), .Q(n8892) );
  HS65_LL_DFPQX4 clk_r_REG98_S2 ( .D(n8459), .CP(clk), .Q(n8891) );
  HS65_LL_DFPQX4 clk_r_REG102_S2 ( .D(n8460), .CP(clk), .Q(n8890) );
  HS65_LL_DFPQX4 clk_r_REG89_S3 ( .D(n8470), .CP(clk), .Q(n8889) );
  HS65_LL_DFPQX4 clk_r_REG70_S2 ( .D(n8472), .CP(clk), .Q(n8888) );
  HS65_LL_DFPQX4 clk_r_REG55_S3 ( .D(n8468), .CP(clk), .Q(n8887) );
  HS65_LL_DFPQX4 clk_r_REG495_S3 ( .D(n8127), .CP(clk), .Q(n8886) );
  HS65_LL_DFPQX4 clk_r_REG494_S3 ( .D(n8080), .CP(clk), .Q(n8885) );
  HS65_LL_DFPQX4 clk_r_REG382_S3 ( .D(n8576), .CP(clk), .Q(n8884) );
  HS65_LL_DFPQNX27 clk_r_REG1_S1 ( .D(\u_DataPath/u_exmemreg/N78 ), .CP(clk), 
        .QN(n7835) );
  HS65_LL_DFPQX4 clk_r_REG35_S2 ( .D(n7839), .CP(clk), .Q(n8883) );
  HS65_LL_DFPQX4 clk_r_REG69_S2 ( .D(n8437), .CP(clk), .Q(n8882) );
  HS65_LL_DFPQX4 clk_r_REG57_S4 ( .D(\lte_x_59/B[5] ), .CP(clk), .Q(n8881) );
  HS65_LL_DFPQX4 clk_r_REG390_S3 ( .D(n8401), .CP(clk), .Q(n8880) );
  HS65_LL_DFPQX4 clk_r_REG294_S1 ( .D(\u_DataPath/mem_writedata_out_i [4]), 
        .CP(clk), .Q(n8879) );
  HS65_LL_DFPQX4 clk_r_REG493_S3 ( .D(n8077), .CP(clk), .Q(n8878) );
  HS65_LL_DFPQX4 clk_r_REG492_S3 ( .D(n8094), .CP(clk), .Q(n8877) );
  HS65_LL_DFPQX4 clk_r_REG50_S1 ( .D(n8428), .CP(clk), .Q(n8875) );
  HS65_LL_DFPQX4 clk_r_REG290_S2 ( .D(\u_DataPath/mem_writedata_out_i [19]), 
        .CP(clk), .Q(n8874) );
  HS65_LL_DFPQX4 clk_r_REG398_S2 ( .D(\u_DataPath/mem_writedata_out_i [2]), 
        .CP(clk), .Q(n8873) );
  HS65_LL_DFPQX4 clk_r_REG295_S2 ( .D(\lte_x_59/B[4] ), .CP(clk), .Q(n8872) );
  HS65_LL_DFPQX4 clk_r_REG475_S3 ( .D(n8100), .CP(clk), .Q(n8871) );
  HS65_LL_DFPQX4 clk_r_REG147_S2 ( .D(\u_DataPath/u_execute/link_value_i [30]), 
        .CP(clk), .Q(n8869) );
  HS65_LL_DFPQX4 clk_r_REG487_S1 ( .D(n8450), .CP(clk), .Q(n8868) );
  HS65_LL_DFPQX4 clk_r_REG332_S1 ( .D(\u_DataPath/data_read_ex_1_i [4]), .CP(
        clk), .Q(n8867) );
  HS65_LL_DFPQX4 clk_r_REG336_S1 ( .D(\u_DataPath/data_read_ex_2_i [22]), .CP(
        clk), .Q(n8866) );
  HS65_LL_DFPQX4 clk_r_REG349_S1 ( .D(\u_DataPath/data_read_ex_2_i [13]), .CP(
        clk), .Q(n8865) );
  HS65_LL_DFPQX4 clk_r_REG401_S1 ( .D(\u_DataPath/data_read_ex_2_i [11]), .CP(
        clk), .Q(n8864) );
  HS65_LL_DFPQX4 clk_r_REG274_S1 ( .D(\u_DataPath/data_read_ex_2_i [9]), .CP(
        clk), .Q(n8863) );
  HS65_LL_DFPQX4 clk_r_REG51_S1 ( .D(\u_DataPath/data_read_ex_1_i [1]), .CP(
        clk), .Q(n8861) );
  HS65_LL_DFPQX4 clk_r_REG404_S1 ( .D(\u_DataPath/data_read_ex_1_i [8]), .CP(
        clk), .Q(n8860) );
  HS65_LL_DFPQX4 clk_r_REG280_S1 ( .D(\u_DataPath/data_read_ex_1_i [26]), .CP(
        clk), .Q(n8859) );
  HS65_LL_DFPQX4 clk_r_REG439_S1 ( .D(\u_DataPath/data_read_ex_1_i [3]), .CP(
        clk), .Q(n8858) );
  HS65_LL_DFPQX4 clk_r_REG360_S1 ( .D(\u_DataPath/data_read_ex_1_i [6]), .CP(
        clk), .Q(n8857) );
  HS65_LL_DFPQX4 clk_r_REG422_S1 ( .D(\u_DataPath/data_read_ex_1_i [12]), .CP(
        clk), .Q(n8856) );
  HS65_LL_DFPQX4 clk_r_REG424_S1 ( .D(\u_DataPath/data_read_ex_1_i [7]), .CP(
        clk), .Q(n8855) );
  HS65_LL_DFPQX4 clk_r_REG288_S1 ( .D(\u_DataPath/data_read_ex_1_i [19]), .CP(
        clk), .Q(n8854) );
  HS65_LL_DFPQX4 clk_r_REG14_S2 ( .D(n8476), .CP(clk), .Q(n8853) );
  HS65_LL_DFPQX4 clk_r_REG11_S3 ( .D(n8467), .CP(clk), .Q(n8852) );
  HS65_LL_DFPQX4 clk_r_REG420_S1 ( .D(\u_DataPath/data_read_ex_1_i [14]), .CP(
        clk), .Q(n8851) );
  HS65_LL_DFPQX4 clk_r_REG348_S1 ( .D(\u_DataPath/data_read_ex_1_i [13]), .CP(
        clk), .Q(n8850) );
  HS65_LL_DFPQX4 clk_r_REG423_S1 ( .D(\u_DataPath/data_read_ex_2_i [12]), .CP(
        clk), .Q(n8849) );
  HS65_LL_DFPQX4 clk_r_REG362_S1 ( .D(\u_DataPath/data_read_ex_2_i [5]), .CP(
        clk), .Q(n8847) );
  HS65_LL_DFPQX4 clk_r_REG342_S1 ( .D(\u_DataPath/data_read_ex_1_i [24]), .CP(
        clk), .Q(n8846) );
  HS65_LL_DFPQX4 clk_r_REG335_S1 ( .D(\u_DataPath/data_read_ex_1_i [22]), .CP(
        clk), .Q(n8845) );
  HS65_LL_DFPQX4 clk_r_REG426_S1 ( .D(\u_DataPath/data_read_ex_2_i [7]), .CP(
        clk), .Q(n8844) );
  HS65_LL_DFPQX4 clk_r_REG414_S1 ( .D(\u_DataPath/data_read_ex_2_i [18]), .CP(
        clk), .Q(n8843) );
  HS65_LL_DFPQX4 clk_r_REG289_S1 ( .D(\u_DataPath/data_read_ex_2_i [19]), .CP(
        clk), .Q(n8842) );
  HS65_LL_DFPQX4 clk_r_REG411_S1 ( .D(\u_DataPath/data_read_ex_1_i [27]), .CP(
        clk), .Q(n8841) );
  HS65_LL_DFPQX4 clk_r_REG380_S1 ( .D(\u_DataPath/data_read_ex_2_i [1]), .CP(
        clk), .Q(n8840) );
  HS65_LL_DFPQX4 clk_r_REG281_S1 ( .D(\u_DataPath/data_read_ex_2_i [23]), .CP(
        clk), .Q(n8839) );
  HS65_LL_DFPQX4 clk_r_REG416_S1 ( .D(\u_DataPath/data_read_ex_1_i [16]), .CP(
        clk), .Q(n8838) );
  HS65_LL_DFPQX4 clk_r_REG291_S1 ( .D(\u_DataPath/data_read_ex_2_i [17]), .CP(
        clk), .Q(n8837) );
  HS65_LL_DFPQX4 clk_r_REG276_S1 ( .D(\u_DataPath/data_read_ex_1_i [21]), .CP(
        clk), .Q(n8836) );
  HS65_LL_DFPQX4 clk_r_REG359_S1 ( .D(\u_DataPath/data_read_ex_2_i [6]), .CP(
        clk), .Q(n8835) );
  HS65_LL_DFPQX4 clk_r_REG338_S1 ( .D(\u_DataPath/data_read_ex_2_i [25]), .CP(
        clk), .Q(n8833) );
  HS65_LL_DFPQX4 clk_r_REG397_S1 ( .D(\u_DataPath/data_read_ex_2_i [31]), .CP(
        clk), .Q(n8832) );
  HS65_LL_DFPQX4 clk_r_REG37_S1 ( .D(\u_DataPath/data_read_ex_1_i [11]), .CP(
        clk), .Q(n8831) );
  HS65_LL_DFPQX4 clk_r_REG405_S1 ( .D(\u_DataPath/data_read_ex_2_i [8]), .CP(
        clk), .Q(n8830) );
  HS65_LL_DFPQX4 clk_r_REG488_S3 ( .D(n8087), .CP(clk), .Q(n8829) );
  HS65_LL_DFPQX4 clk_r_REG54_S3 ( .D(n7848), .CP(clk), .Q(n8828) );
  HS65_LL_DFPRQX4 clk_r_REG192_S5 ( .D(\u_DataPath/pc4_to_idexreg_i [31]), 
        .CP(clk), .RN(n8676), .Q(n8827) );
  HS65_LL_DFPQX4 clk_r_REG67_S1 ( .D(\u_DataPath/data_read_ex_1_i [29]), .CP(
        clk), .Q(n8826) );
  HS65_LL_DFPQX4 clk_r_REG286_S1 ( .D(\u_DataPath/data_read_ex_1_i [20]), .CP(
        clk), .Q(n8825) );
  HS65_LL_DFPQX4 clk_r_REG413_S1 ( .D(\u_DataPath/data_read_ex_1_i [18]), .CP(
        clk), .Q(n8824) );
  HS65_LL_DFPQX4 clk_r_REG396_S1 ( .D(\u_DataPath/data_read_ex_1_i [31]), .CP(
        clk), .Q(n8823) );
  HS65_LL_DFPQX4 clk_r_REG91_S1 ( .D(\u_DataPath/data_read_ex_1_i [17]), .CP(
        clk), .Q(n8822) );
  HS65_LL_DFPQX4 clk_r_REG357_S2 ( .D(\u_DataPath/data_read_ex_1_i [28]), .CP(
        clk), .Q(n8821) );
  HS65_LL_DFPRQX4 clk_r_REG610_S3 ( .D(\u_DataPath/immediate_ext_dec_i [15]), 
        .CP(clk), .RN(n9354), .Q(n8818) );
  HS65_LL_DFPRQX4 clk_r_REG131_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [14]), 
        .CP(clk), .RN(n8676), .Q(n8815) );
  HS65_LL_DFPRQX4 clk_r_REG250_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [15]), 
        .CP(clk), .RN(n9361), .Q(n8814) );
  HS65_LL_DFPRQX4 clk_r_REG372_S3 ( .D(\u_DataPath/pc4_to_idexreg_i [2]), .CP(
        clk), .RN(n2877), .Q(n8811) );
  HS65_LL_DFPRQX4 clk_r_REG4_S3 ( .D(\u_DataPath/pc4_to_idexreg_i [3]), .CP(
        clk), .RN(n9361), .Q(n8810) );
  HS65_LL_DFPQX4 clk_r_REG88_S3 ( .D(n8462), .CP(clk), .Q(n8801) );
  HS65_LL_DFPQX4 clk_r_REG273_S1 ( .D(\u_DataPath/data_read_ex_1_i [9]), .CP(
        clk), .Q(n8800) );
  HS65_LL_DFPQX4 clk_r_REG84_S1 ( .D(\u_DataPath/data_read_ex_1_i [25]), .CP(
        clk), .Q(n8799) );
  HS65_LL_DFPQX4 clk_r_REG400_S1 ( .D(\u_DataPath/data_read_ex_1_i [2]), .CP(
        clk), .Q(n8798) );
  HS65_LL_DFPRQX4 clk_r_REG199_S5 ( .D(\u_DataPath/pc4_to_idexreg_i [29]), 
        .CP(clk), .RN(n9361), .Q(n8796) );
  HS65_LL_DFPRQX4 clk_r_REG236_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [17]), 
        .CP(clk), .RN(n8676), .Q(n8795) );
  HS65_LL_DFPQX4 clk_r_REG526_S2 ( .D(opcode_i[3]), .CP(clk), .Q(n8794) );
  HS65_LL_DFPRQX4 clk_r_REG607_S3 ( .D(\u_DataPath/immediate_ext_dec_i [14]), 
        .CP(clk), .RN(n9354), .Q(n8791) );
  HS65_LL_DFPRQX4 clk_r_REG601_S3 ( .D(\u_DataPath/immediate_ext_dec_i [12]), 
        .CP(clk), .RN(n9354), .Q(n8789) );
  HS65_LL_DFPRQX4 clk_r_REG598_S3 ( .D(\u_DataPath/immediate_ext_dec_i [11]), 
        .CP(clk), .RN(n9354), .Q(n8788) );
  HS65_LL_DFPRQX4 clk_r_REG595_S3 ( .D(\u_DataPath/immediate_ext_dec_i [4]), 
        .CP(clk), .RN(n9354), .Q(n8780) );
  HS65_LL_DFPRQX4 clk_r_REG590_S3 ( .D(\u_DataPath/immediate_ext_dec_i [5]), 
        .CP(clk), .RN(n9354), .Q(n8779) );
  HS65_LL_DFPRQX4 clk_r_REG587_S3 ( .D(\u_DataPath/immediate_ext_dec_i [6]), 
        .CP(clk), .RN(n9354), .Q(n8778) );
  HS65_LL_DFPQX4 clk_r_REG584_S3 ( .D(\u_DataPath/immediate_ext_dec_i [0]), 
        .CP(clk), .Q(n8777) );
  HS65_LL_DFPRQX4 clk_r_REG583_S3 ( .D(\u_DataPath/immediate_ext_dec_i [0]), 
        .CP(clk), .RN(n9354), .Q(n8776) );
  HS65_LL_DFPQX4 clk_r_REG577_S3 ( .D(\u_DataPath/immediate_ext_dec_i [1]), 
        .CP(clk), .Q(n8775) );
  HS65_LL_DFPRQX4 clk_r_REG576_S3 ( .D(\u_DataPath/immediate_ext_dec_i [1]), 
        .CP(clk), .RN(n9354), .Q(n8774) );
  HS65_LL_DFPRQX4 clk_r_REG569_S3 ( .D(\u_DataPath/immediate_ext_dec_i [3]), 
        .CP(clk), .RN(n9354), .Q(n8772) );
  HS65_LL_DFPQX4 clk_r_REG564_S3 ( .D(\u_DataPath/immediate_ext_dec_i [2]), 
        .CP(clk), .Q(n8771) );
  HS65_LL_DFPRQX4 clk_r_REG563_S3 ( .D(\u_DataPath/immediate_ext_dec_i [2]), 
        .CP(clk), .RN(n9354), .Q(n8770) );
  HS65_LL_DFPQX4 clk_r_REG491_S3 ( .D(n8099), .CP(clk), .Q(n8767) );
  HS65_LL_DFPQX4 clk_r_REG504_S1 ( .D(\u_DataPath/RFaddr_out_memwb_i [1]), 
        .CP(clk), .Q(n8766) );
  HS65_LL_DFPQX4 clk_r_REG502_S1 ( .D(\u_DataPath/RFaddr_out_memwb_i [2]), 
        .CP(clk), .Q(n8764) );
  HS65_LL_DFPQX4 clk_r_REG500_S1 ( .D(\u_DataPath/RFaddr_out_memwb_i [0]), 
        .CP(clk), .Q(n8763) );
  HS65_LL_DFPQX4 clk_r_REG498_S1 ( .D(\u_DataPath/RFaddr_out_memwb_i [4]), 
        .CP(clk), .Q(n8762) );
  HS65_LL_DFPQX4 clk_r_REG496_S1 ( .D(\u_DataPath/RFaddr_out_memwb_i [3]), 
        .CP(clk), .Q(n8761) );
  HS65_LL_DFPQX4 clk_r_REG78_S2 ( .D(n8309), .CP(clk), .Q(n8760) );
  HS65_LL_DFPQX4 clk_r_REG352_S2 ( .D(n8296), .CP(clk), .Q(n8759) );
  HS65_LL_DFPQX4 clk_r_REG386_S2 ( .D(n8169), .CP(clk), .Q(n8758) );
  HS65_LL_DFPRQX4 clk_r_REG561_S3 ( .D(\u_DataPath/jaddr_i [25]), .CP(clk), 
        .RN(n9354), .Q(n8756) );
  HS65_LL_DFPQX4 clk_r_REG486_S3 ( .D(\u_DataPath/cw_to_ex_i [17]), .CP(clk), 
        .Q(n8755) );
  HS65_LL_DFPRQX4 clk_r_REG533_S2 ( .D(\u_DataPath/jaddr_i [16]), .CP(clk), 
        .RN(n9354), .Q(n8754) );
  HS65_LL_DFPQX4 clk_r_REG351_S2 ( .D(n8181), .CP(clk), .Q(n8753) );
  HS65_LL_DFPQX4 clk_r_REG344_S2 ( .D(n8305), .CP(clk), .Q(n8752) );
  HS65_LL_DFPQX4 clk_r_REG481_S3 ( .D(n8057), .CP(clk), .Q(n8750) );
  HS65_LL_DFPQX4 clk_r_REG65_S2 ( .D(\u_DataPath/mem_writedata_out_i [29]), 
        .CP(clk), .Q(n8749) );
  HS65_LL_DFPQX4 clk_r_REG285_S2 ( .D(\u_DataPath/mem_writedata_out_i [20]), 
        .CP(clk), .Q(n8747) );
  HS65_LL_DFPQX4 clk_r_REG106_S2 ( .D(\u_DataPath/mem_writedata_out_i [21]), 
        .CP(clk), .Q(n8746) );
  HS65_LL_DFPQX4 clk_r_REG13_S2 ( .D(\u_DataPath/mem_writedata_out_i [7]), 
        .CP(clk), .Q(n8745) );
  HS65_LL_DFPQX4 clk_r_REG381_S2 ( .D(\u_DataPath/mem_writedata_out_i [1]), 
        .CP(clk), .Q(n8744) );
  HS65_LL_DFPQX4 clk_r_REG358_S2 ( .D(\u_DataPath/mem_writedata_out_i [6]), 
        .CP(clk), .Q(n8743) );
  HS65_LL_DFPQX4 clk_r_REG75_S1 ( .D(\u_DataPath/mem_writedata_out_i [13]), 
        .CP(clk), .Q(n8742) );
  HS65_LL_DFPQX4 clk_r_REG72_S1 ( .D(\u_DataPath/mem_writedata_out_i [10]), 
        .CP(clk), .Q(n8741) );
  HS65_LL_DFPQX4 clk_r_REG418_S1 ( .D(\u_DataPath/mem_writedata_out_i [14]), 
        .CP(clk), .Q(n8739) );
  HS65_LL_DFPQX4 clk_r_REG23_S1 ( .D(\u_DataPath/mem_writedata_out_i [16]), 
        .CP(clk), .Q(n8738) );
  HS65_LL_DFPQX4 clk_r_REG415_S1 ( .D(\u_DataPath/mem_writedata_out_i [18]), 
        .CP(clk), .Q(n8737) );
  HS65_LL_DFPQX4 clk_r_REG282_S1 ( .D(\u_DataPath/mem_writedata_out_i [23]), 
        .CP(clk), .Q(n8736) );
  HS65_LL_DFPQX4 clk_r_REG402_S1 ( .D(\u_DataPath/mem_writedata_out_i [11]), 
        .CP(clk), .Q(n8735) );
  HS65_LL_DFPQX4 clk_r_REG345_S1 ( .D(\u_DataPath/mem_writedata_out_i [15]), 
        .CP(clk), .Q(n8734) );
  HS65_LL_DFPQX4 clk_r_REG278_S1 ( .D(\u_DataPath/mem_writedata_out_i [26]), 
        .CP(clk), .Q(n8733) );
  HS65_LL_DFPQX4 clk_r_REG363_S1 ( .D(\u_DataPath/mem_writedata_out_i [5]), 
        .CP(clk), .Q(n8731) );
  HS65_LL_DFPQX4 clk_r_REG16_S1 ( .D(\u_DataPath/mem_writedata_out_i [12]), 
        .CP(clk), .Q(n8730) );
  HS65_LL_DFPQX4 clk_r_REG408_S1 ( .D(\u_DataPath/mem_writedata_out_i [30]), 
        .CP(clk), .Q(n8729) );
  HS65_LL_DFPQX4 clk_r_REG44_S1 ( .D(\u_DataPath/mem_writedata_out_i [31]), 
        .CP(clk), .Q(n8728) );
  HS65_LL_DFPQX4 clk_r_REG334_S1 ( .D(\u_DataPath/mem_writedata_out_i [22]), 
        .CP(clk), .Q(n8727) );
  HS65_LL_DFPQX4 clk_r_REG272_S1 ( .D(\u_DataPath/mem_writedata_out_i [9]), 
        .CP(clk), .Q(n8726) );
  HS65_LL_DFPQX4 clk_r_REG331_S1 ( .D(\u_DataPath/data_read_ex_2_i [4]), .CP(
        clk), .Q(n8724) );
  HS65_LL_DFPQX4 clk_r_REG419_S1 ( .D(\u_DataPath/data_read_ex_2_i [14]), .CP(
        clk), .Q(n8723) );
  HS65_LL_DFPQX4 clk_r_REG407_S1 ( .D(\u_DataPath/data_read_ex_2_i [30]), .CP(
        clk), .Q(n8722) );
  HS65_LL_DFPQX4 clk_r_REG410_S1 ( .D(\u_DataPath/data_read_ex_2_i [27]), .CP(
        clk), .Q(n8721) );
  HS65_LL_DFPQX4 clk_r_REG284_S1 ( .D(\u_DataPath/data_read_ex_2_i [20]), .CP(
        clk), .Q(n8720) );
  HS65_LL_DFPQX4 clk_r_REG66_S1 ( .D(\u_DataPath/data_read_ex_2_i [29]), .CP(
        clk), .Q(n8719) );
  HS65_LL_DFPQX4 clk_r_REG22_S1 ( .D(\u_DataPath/data_read_ex_2_i [16]), .CP(
        clk), .Q(n8718) );
  HS65_LL_DFPQX4 clk_r_REG275_S1 ( .D(\u_DataPath/data_read_ex_2_i [21]), .CP(
        clk), .Q(n8717) );
  HS65_LL_DFPQX4 clk_r_REG399_S1 ( .D(\u_DataPath/data_read_ex_2_i [2]), .CP(
        clk), .Q(n8716) );
  HS65_LL_DFPQX4 clk_r_REG49_S1 ( .D(\u_DataPath/u_execute/psw_status_i [0]), 
        .CP(clk), .Q(n8715) );
  HS65_LL_DFPQX4 clk_r_REG480_S3 ( .D(n8102), .CP(clk), .Q(n8702) );
  HS65_LL_DFPQX4 clk_r_REG474_S3 ( .D(n8081), .CP(clk), .Q(n8696) );
  HS65_LH_IVX2 U3797 ( .A(n9330), .Z(n8676) );
  HS65_LH_IVX2 U3799 ( .A(n9330), .Z(n8677) );
  HS65_LH_IVX2 U5114 ( .A(n2877), .Z(n9330) );
  HS65_LH_DFPHQX4 clk_r_REG190_S3 ( .D(n8641), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8713) );
  HS65_LH_DFPRQX4 clk_r_REG537_S2 ( .D(n8482), .CP(clk), .RN(n9356), .Q(n9069)
         );
  HS65_LH_DFPRQX4 clk_r_REG428_S2 ( .D(n8691), .CP(clk), .RN(n8676), .Q(n8690)
         );
  HS65_LH_DFPRQX4 clk_r_REG365_S2 ( .D(n8689), .CP(clk), .RN(n9361), .Q(n8688)
         );
  HS65_LH_DFPRQX4 clk_r_REG646_S1 ( .D(iram_data[0]), .CP(clk), .RN(n9355), 
        .Q(n9303) );
  HS65_LH_DFPRQX4 clk_r_REG645_S1 ( .D(iram_data[1]), .CP(clk), .RN(n9356), 
        .Q(n9304) );
  HS65_LH_DFPRQX4 clk_r_REG644_S1 ( .D(iram_data[2]), .CP(clk), .RN(n9355), 
        .Q(n9305) );
  HS65_LH_DFPRQX4 clk_r_REG643_S1 ( .D(iram_data[3]), .CP(clk), .RN(n9356), 
        .Q(n9306) );
  HS65_LH_DFPRQX4 clk_r_REG642_S1 ( .D(iram_data[4]), .CP(clk), .RN(n9355), 
        .Q(n9307) );
  HS65_LH_DFPRQX4 clk_r_REG641_S1 ( .D(iram_data[5]), .CP(clk), .RN(n9356), 
        .Q(n9308) );
  HS65_LH_DFPRQX4 clk_r_REG640_S1 ( .D(iram_data[6]), .CP(clk), .RN(n9355), 
        .Q(n9309) );
  HS65_LH_DFPRQX4 clk_r_REG638_S1 ( .D(iram_data[8]), .CP(clk), .RN(n9354), 
        .Q(n9311) );
  HS65_LH_DFPRQX4 clk_r_REG637_S1 ( .D(iram_data[9]), .CP(clk), .RN(n9361), 
        .Q(n9312) );
  HS65_LH_DFPRQX4 clk_r_REG635_S1 ( .D(iram_data[11]), .CP(clk), .RN(n9356), 
        .Q(n9314) );
  HS65_LH_DFPRQX4 clk_r_REG634_S1 ( .D(iram_data[12]), .CP(clk), .RN(n9355), 
        .Q(n9315) );
  HS65_LH_DFPRQX4 clk_r_REG633_S1 ( .D(iram_data[13]), .CP(clk), .RN(n9356), 
        .Q(n9316) );
  HS65_LH_DFPRQX4 clk_r_REG632_S1 ( .D(iram_data[14]), .CP(clk), .RN(n9355), 
        .Q(n9317) );
  HS65_LH_DFPRQX4 clk_r_REG631_S1 ( .D(iram_data[15]), .CP(clk), .RN(n9356), 
        .Q(n9318) );
  HS65_LH_DFPRQX4 clk_r_REG630_S1 ( .D(iram_data[16]), .CP(clk), .RN(n9355), 
        .Q(n9319) );
  HS65_LH_DFPRQX4 clk_r_REG629_S1 ( .D(iram_data[17]), .CP(clk), .RN(n9356), 
        .Q(n9320) );
  HS65_LH_DFPRQX4 clk_r_REG628_S1 ( .D(iram_data[18]), .CP(clk), .RN(n9355), 
        .Q(n9321) );
  HS65_LH_DFPRQX4 clk_r_REG627_S1 ( .D(iram_data[19]), .CP(clk), .RN(n9356), 
        .Q(n9322) );
  HS65_LH_DFPRQX4 clk_r_REG626_S1 ( .D(iram_data[20]), .CP(clk), .RN(n9355), 
        .Q(n9323) );
  HS65_LH_DFPRQX4 clk_r_REG625_S1 ( .D(iram_data[21]), .CP(clk), .RN(n9356), 
        .Q(n9324) );
  HS65_LH_DFPRQX4 clk_r_REG624_S1 ( .D(iram_data[22]), .CP(clk), .RN(n9355), 
        .Q(n9325) );
  HS65_LH_DFPRQX4 clk_r_REG623_S1 ( .D(iram_data[23]), .CP(clk), .RN(n9356), 
        .Q(n9326) );
  HS65_LH_DFPRQX4 clk_r_REG622_S1 ( .D(iram_data[24]), .CP(clk), .RN(n9355), 
        .Q(n9327) );
  HS65_LH_DFPRQX4 clk_r_REG621_S1 ( .D(iram_data[25]), .CP(clk), .RN(n9356), 
        .Q(n9328) );
  HS65_LH_DFPRQX4 clk_r_REG620_S1 ( .D(iram_data[27]), .CP(clk), .RN(n9355), 
        .Q(n9329) );
  HS65_LH_DFPRQX4 clk_r_REG619_S1 ( .D(iram_data[29]), .CP(clk), .RN(n9356), 
        .Q(n9331) );
  HS65_LH_DFPRQX4 clk_r_REG544_S3 ( .D(\u_DataPath/immediate_ext_dec_i [8]), 
        .CP(clk), .RN(n8676), .Q(n8783) );
  HS65_LH_DFPRQX4 clk_r_REG547_S3 ( .D(\u_DataPath/immediate_ext_dec_i [9]), 
        .CP(clk), .RN(n9361), .Q(n8782) );
  HS65_LH_DFPRQX4 clk_r_REG155_S5 ( .D(n9429), .CP(clk), .RN(n9355), .Q(n9159)
         );
  HS65_LH_DFPRQX4 clk_r_REG138_S4 ( .D(n9428), .CP(clk), .RN(n9356), .Q(n9163)
         );
  HS65_LH_DFPRQX4 clk_r_REG516_S2 ( .D(opcode_i[5]), .CP(clk), .RN(n8676), .Q(
        n8786) );
  HS65_LH_DFPRQX4 clk_r_REG265_S4 ( .D(n9422), .CP(clk), .RN(n9361), .Q(n9158)
         );
  HS65_LH_DFPRQX4 clk_r_REG215_S4 ( .D(n9426), .CP(clk), .RN(n8676), .Q(n9156)
         );
  HS65_LH_DFPRQX4 clk_r_REG208_S5 ( .D(n9420), .CP(clk), .RN(n9361), .Q(n9161)
         );
  HS65_LH_DFPRQX4 clk_r_REG170_S5 ( .D(n9427), .CP(clk), .RN(n8676), .Q(n9155)
         );
  HS65_LH_DFPRQX4 clk_r_REG113_S5 ( .D(n9423), .CP(clk), .RN(n9361), .Q(n9157)
         );
  HS65_LH_DFPRQX4 clk_r_REG519_S2 ( .D(\u_DataPath/jaddr_i [23]), .CP(clk), 
        .RN(n9355), .Q(n8820) );
  HS65_LH_DFPRQX4 clk_r_REG525_S2 ( .D(opcode_i[3]), .CP(clk), .RN(n9355), .Q(
        n8793) );
  HS65_LH_DFPRQX4 clk_r_REG528_S2 ( .D(opcode_i[1]), .CP(clk), .RN(n9356), .Q(
        n8792) );
  HS65_LH_DFPRQX4 clk_r_REG521_S2 ( .D(\u_DataPath/jaddr_i [21]), .CP(clk), 
        .RN(n9356), .Q(n8817) );
  HS65_LH_DFPRQX4 clk_r_REG557_S3 ( .D(\u_DataPath/jaddr_i [24]), .CP(clk), 
        .RN(n9355), .Q(n8819) );
  HS65_LH_DFPRQX4 clk_r_REG553_S3 ( .D(\u_DataPath/jaddr_i [18]), .CP(clk), 
        .RN(n9356), .Q(n8787) );
  HS65_LH_DFPRQX4 clk_r_REG523_S2 ( .D(\u_DataPath/jaddr_i [20]), .CP(clk), 
        .RN(n9355), .Q(n8816) );
  HS65_LH_DFPRQX4 clk_r_REG297_S4 ( .D(\u_DataPath/pc_4_i [4]), .CP(clk), .RN(
        n8676), .Q(n9009) );
  HS65_LH_DFPRQX4 clk_r_REG529_S2 ( .D(\u_DataPath/jaddr_i [19]), .CP(clk), 
        .RN(n9356), .Q(n8785) );
  HS65_LH_DFPRQX4 clk_r_REG531_S2 ( .D(\u_DataPath/jaddr_i [17]), .CP(clk), 
        .RN(n9355), .Q(n8757) );
  HS65_LH_DFPRQX4 clk_r_REG326_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [5]), .CP(
        clk), .RN(n9361), .Q(n8809) );
  HS65_LH_DFPRQX4 clk_r_REG307_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [6]), .CP(
        clk), .RN(n8676), .Q(n8807) );
  HS65_LH_DFPRQX4 clk_r_REG298_S5 ( .D(\u_DataPath/pc4_to_idexreg_i [4]), .CP(
        clk), .RN(n9361), .Q(n8768) );
  HS65_LH_DFPSQX4 clk_r_REG507_S2 ( .D(opcode_i[0]), .CP(clk), .SN(n7879), .Q(
        n9084) );
  HS65_LH_DFPSQX4 clk_r_REG455_S2 ( .D(opcode_i[2]), .CP(clk), .SN(n7879), .Q(
        n9082) );
  HS65_LH_DFPSQX4 clk_r_REG440_S2 ( .D(opcode_i[4]), .CP(clk), .SN(n7879), .Q(
        n9068) );
  HS65_LH_DFPHQX4 clk_r_REG427_S1 ( .D(\u_DataPath/pc_4_i [0]), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n8691) );
  HS65_LH_DFPHQX4 clk_r_REG370_S1 ( .D(n8670), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8687) );
  HS65_LH_DFPHQX4 clk_r_REG364_S1 ( .D(\u_DataPath/pc_4_i [1]), .E(
        \u_DataPath/u_fetch/pc1/N3 ), .CP(clk), .Q(n8689) );
  HS65_LH_DFPHQX4 clk_r_REG324_S2 ( .D(n8667), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8684) );
  HS65_LH_DFPHQX4 clk_r_REG316_S2 ( .D(n8665), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8682) );
  HS65_LH_DFPHQX4 clk_r_REG310_S2 ( .D(n8664), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8680) );
  HS65_LH_DFPHQX4 clk_r_REG305_S2 ( .D(n8666), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8683) );
  HS65_LH_DFPHQX4 clk_r_REG296_S3 ( .D(n8668), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8685) );
  HS65_LH_DFPHQX4 clk_r_REG263_S2 ( .D(n8661), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8679) );
  HS65_LH_DFPHQX4 clk_r_REG117_S2 ( .D(n8662), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8681) );
  HS65_LH_DFPHQX4 clk_r_REG111_S3 ( .D(n8663), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8678) );
  HS65_LH_DFPHQX4 clk_r_REG2_S1 ( .D(n8669), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8686) );
  HS65_LH_DFPHQX4 clk_r_REG256_S2 ( .D(n8660), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8695) );
  HS65_LH_DFPHQX4 clk_r_REG129_S2 ( .D(n8658), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8694) );
  HS65_LH_DFPHQX4 clk_r_REG123_S2 ( .D(n8659), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8698) );
  HS65_LH_DFPHQX4 clk_r_REG213_S2 ( .D(n8654), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8693) );
  HS65_LH_DFPHQX4 clk_r_REG168_S3 ( .D(n8646), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8701) );
  HS65_LH_DFPHQX4 clk_r_REG248_S2 ( .D(n8657), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8699) );
  HS65_LH_DFPHQX4 clk_r_REG174_S2 ( .D(n8645), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8703) );
  HS65_LH_DFPHQX4 clk_r_REG241_S2 ( .D(n8656), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8704) );
  HS65_LH_DFPHQX4 clk_r_REG221_S2 ( .D(n8653), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8692) );
  HS65_LH_DFPHQX4 clk_r_REG163_S3 ( .D(n8647), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8700) );
  HS65_LH_DFPHQX4 clk_r_REG226_S2 ( .D(n8652), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8697) );
  HS65_LH_DFPHQX4 clk_r_REG180_S3 ( .D(n8644), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8707) );
  HS65_LH_DFPHQX4 clk_r_REG234_S2 ( .D(n8655), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8709) );
  HS65_LH_DFPHQX4 clk_r_REG153_S3 ( .D(n8650), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8708) );
  HS65_LH_DFPHQX4 clk_r_REG197_S3 ( .D(n8643), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8710) );
  HS65_LH_DFPHQX4 clk_r_REG206_S3 ( .D(n8649), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8706) );
  HS65_LH_DFPHQX4 clk_r_REG158_S3 ( .D(n8648), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8711) );
  HS65_LH_DFPHQX4 clk_r_REG185_S3 ( .D(n8642), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8712) );
  HS65_LH_DFPHQX4 clk_r_REG136_S2 ( .D(n8651), .E(\u_DataPath/u_fetch/pc1/N3 ), 
        .CP(clk), .Q(n8705) );
  HS65_LH_DFPQX4 clk_r_REG46_S2 ( .D(n9118), .CP(clk), .Q(n9117) );
  HS65_LL_DFPQNX4 clk_r_REG466_S1 ( .D(n8048), .CP(clk), .QN(
        \u_DataPath/cw_towb_i [1]) );
  HS65_LH_DFPQX9 clk_r_REG436_S3 ( .D(nibble[0]), .CP(clk), .Q(n9128) );
  HS65_LL_DFPRQX9 clk_r_REG613_S1 ( .D(n7923), .CP(clk), .RN(n9356), .Q(n9252)
         );
  HS65_LL_DFPQX9 clk_r_REG562_S1 ( .D(n8626), .CP(clk), .Q(n8911) );
  HS65_LH_DFPQX9 clk_r_REG541_S3 ( .D(n8073), .CP(clk), .Q(n8751) );
  HS65_LH_DFPQX9 clk_r_REG591_S3 ( .D(n8074), .CP(clk), .Q(n9002) );
  HS65_LH_DFPQX9 clk_r_REG582_S3 ( .D(n8123), .CP(clk), .Q(n9146) );
  HS65_LH_DFPQX9 clk_r_REG482_S4 ( .D(\u_DataPath/u_idexreg/N184 ), .CP(clk), 
        .Q(n8876) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][12]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7968), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][12] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][8]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7939), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][28]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7929), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][28] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][7]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7950), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][7] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7956), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][30]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n8012), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][30] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][20]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7959), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][20] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7983), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][13]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7957), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][13] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7989), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][14] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][14]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7990), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ) );
  HS65_LH_DFPQX4 clk_r_REG665_S1 ( .D(Data_out_fromRAM[21]), .CP(clk), .Q(
        n9294) );
  HS65_LH_DFPQX4 clk_r_REG687_S1 ( .D(Data_out_fromRAM[5]), .CP(clk), .Q(n9279) );
  HS65_LH_DFPQX4 clk_r_REG287_S3 ( .D(n2849), .CP(clk), .Q(n9262) );
  HS65_LH_DFPQX4 clk_r_REG653_S1 ( .D(n8417), .CP(clk), .Q(n9246) );
  HS65_LH_DFPQX4 clk_r_REG114_S1 ( .D(\u_DataPath/pc_4_to_ex_i [9]), .CP(clk), 
        .Q(n9231) );
  HS65_LH_DFPQX4 clk_r_REG139_S1 ( .D(\u_DataPath/pc_4_to_ex_i [21]), .CP(clk), 
        .Q(n9216) );
  HS65_LH_DFPQX4 clk_r_REG101_S3 ( .D(n7838), .CP(clk), .Q(n9201) );
  HS65_LH_DFPQX4 clk_r_REG353_S1 ( .D(n7947), .CP(clk), .Q(n9186) );
  HS65_LH_DFPQX4 clk_r_REG551_S1 ( .D(\u_DataPath/immediate_ext_ex_i [10]), 
        .CP(clk), .Q(n9171) );
  HS65_LH_DFPQX4 clk_r_REG377_S1 ( .D(\u_DataPath/branch_target_i [3]), .CP(
        clk), .Q(n9147) );
  HS65_LH_DFPQX4 clk_r_REG617_S1 ( .D(n8058), .CP(clk), .Q(n9130) );
  HS65_LH_DFPQX4 clk_r_REG478_S1 ( .D(\u_DataPath/cw_tomem_i [5]), .CP(clk), 
        .Q(n9113) );
  HS65_LH_DFPRQX9 clk_r_REG317_S3 ( .D(\u_DataPath/pc_4_i [7]), .CP(clk), .RN(
        n9362), .Q(n9098) );
  HS65_LH_DFPQX4 clk_r_REG261_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [12]), 
        .CP(clk), .Q(n9064) );
  HS65_LH_DFPQX4 clk_r_REG585_S1 ( .D(\u_DataPath/immediate_ext_ex_i [0]), 
        .CP(clk), .Q(n9035) );
  HS65_LH_DFPQX4 clk_r_REG150_S2 ( .D(\u_DataPath/u_execute/link_value_i [26]), 
        .CP(clk), .Q(n9020) );
  HS65_LH_DFPRQX4 clk_r_REG112_S4 ( .D(\u_DataPath/pc_4_i [9]), .CP(clk), .RN(
        n2877), .Q(n8973) );
  HS65_LH_DFPQX4 clk_r_REG321_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [6]), 
        .CP(clk), .Q(n8959) );
  HS65_LH_DFPQX4 clk_r_REG211_S1 ( .D(\u_DataPath/branch_target_i [22]), .CP(
        clk), .Q(n8929) );
  HS65_LH_DFPQX4 clk_r_REG485_S1 ( .D(\u_DataPath/cw_tomem_i [3]), .CP(clk), 
        .Q(n8915) );
  HS65_LH_DFPQX4 clk_r_REG59_S1 ( .D(\u_DataPath/from_alu_data_out_i [6]), 
        .CP(clk), .Q(n8908) );
  HS65_LH_DFPQNX4 clk_r_REG28_S1 ( .D(\u_DataPath/from_alu_data_out_i [27]), 
        .CP(clk), .QN(n3020) );
  HS65_LH_DFPQX4 clk_r_REG39_S2 ( .D(n8464), .CP(clk), .Q(n8894) );
  HS65_LH_DFPQX4 clk_r_REG283_S1 ( .D(\u_DataPath/data_read_ex_1_i [23]), .CP(
        clk), .Q(n8848) );
  HS65_LH_DFPQX4 clk_r_REG409_S1 ( .D(\u_DataPath/data_read_ex_1_i [30]), .CP(
        clk), .Q(n8834) );
  HS65_LH_DFPRQX4 clk_r_REG160_S5 ( .D(\u_DataPath/pc4_to_idexreg_i [24]), 
        .CP(clk), .RN(n9361), .Q(n8797) );
  HS65_LH_DFPQX4 clk_r_REG570_S3 ( .D(\u_DataPath/immediate_ext_dec_i [3]), 
        .CP(clk), .Q(n8773) );
  HS65_LH_DFPQX4 clk_r_REG292_S1 ( .D(\u_DataPath/mem_writedata_out_i [17]), 
        .CP(clk), .Q(n8740) );
  HS65_LH_DFPQX4 clk_r_REG438_S1 ( .D(\u_DataPath/mem_writedata_out_i [3]), 
        .CP(clk), .Q(n8725) );
  HS65_LH_DFPQX4 clk_r_REG506_S4 ( .D(\u_DataPath/cw_to_ex_i [15]), .CP(clk), 
        .Q(n8714) );
  HS65_LH_DFPRQX9 clk_r_REG318_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [7]), .CP(
        clk), .RN(n9360), .Q(n8806) );
  HS65_LH_DFPRQX9 clk_r_REG3_S2 ( .D(\u_DataPath/pc_4_i [3]), .CP(clk), .RN(
        n9360), .Q(n8970) );
  HS65_LH_DFPRQX9 clk_r_REG187_S5 ( .D(n9421), .CP(clk), .RN(n9360), .Q(n9143)
         );
  HS65_LH_DFPRQX9 clk_r_REG258_S4 ( .D(n9419), .CP(clk), .RN(n9360), .Q(n9265)
         );
  HS65_LH_DFPRQX9 clk_r_REG550_S3 ( .D(\u_DataPath/immediate_ext_dec_i [10]), 
        .CP(clk), .RN(n9360), .Q(n8781) );
  HS65_LH_DFPRQX9 clk_r_REG371_S2 ( .D(\u_DataPath/pc_4_i [2]), .CP(clk), .RN(
        n9360), .Q(n9273) );
  HS65_LH_DFPRQX9 clk_r_REG223_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [19]), 
        .CP(clk), .RN(n9360), .Q(n8813) );
  HS65_LH_DFPRQX9 clk_r_REG165_S5 ( .D(\u_DataPath/pc4_to_idexreg_i [25]), 
        .CP(clk), .RN(n9360), .Q(n8802) );
  HS65_LH_DFPRQX9 clk_r_REG119_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [10]), 
        .CP(clk), .RN(n9360), .Q(n8804) );
  HS65_LH_DFPRQX9 clk_r_REG325_S3 ( .D(\u_DataPath/pc_4_i [5]), .CP(clk), .RN(
        n9360), .Q(n8971) );
  HS65_LH_DFPRQX9 clk_r_REG311_S3 ( .D(\u_DataPath/pc_4_i [8]), .CP(clk), .RN(
        n9360), .Q(n9010) );
  HS65_LH_DFPRQX9 clk_r_REG130_S3 ( .D(\u_DataPath/pc_4_i [14]), .CP(clk), 
        .RN(n9360), .Q(n8984) );
  HS65_LH_DFPRQX9 clk_r_REG249_S3 ( .D(\u_DataPath/pc_4_i [15]), .CP(clk), 
        .RN(n9360), .Q(n9097) );
  HS65_LH_DFPRQX9 clk_r_REG164_S4 ( .D(\u_DataPath/pc_4_i [25]), .CP(clk), 
        .RN(n9360), .Q(n8980) );
  HS65_LH_DFPRQX9 clk_r_REG198_S4 ( .D(\u_DataPath/pc_4_i [29]), .CP(clk), 
        .RN(n9360), .Q(n8993) );
  HS65_LH_DFPRQX9 clk_r_REG536_S1 ( .D(n7921), .CP(clk), .RN(n9360), .Q(n9192)
         );
  HS65_LH_DFPRQX9 clk_r_REG515_S1 ( .D(n7924), .CP(clk), .RN(n9360), .Q(n9139)
         );
  HS65_LH_DFPRQX9 clk_r_REG556_S2 ( .D(n7918), .CP(clk), .RN(n9360), .Q(n9154)
         );
  HS65_LH_DFPRQX9 clk_r_REG636_S1 ( .D(iram_data[10]), .CP(clk), .RN(n9360), 
        .Q(n9313) );
  HS65_LH_DFPRQX9 clk_r_REG312_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [8]), .CP(
        clk), .RN(n9362), .Q(n8805) );
  HS65_LH_DFPRQX9 clk_r_REG429_S3 ( .D(\u_DataPath/pc4_to_idexreg_i [0]), .CP(
        clk), .RN(n9362), .Q(n8862) );
  HS65_LH_DFPRQX9 clk_r_REG182_S5 ( .D(n9425), .CP(clk), .RN(n9362), .Q(n9160)
         );
  HS65_LH_DFPRQX9 clk_r_REG243_S4 ( .D(n9424), .CP(clk), .RN(n9362), .Q(n9162)
         );
  HS65_LH_DFPRQX9 clk_r_REG540_S3 ( .D(\u_DataPath/immediate_ext_dec_i [7]), 
        .CP(clk), .RN(n9362), .Q(n8784) );
  HS65_LH_DFPRQX9 clk_r_REG228_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [20]), 
        .CP(clk), .RN(n9362), .Q(n8812) );
  HS65_LH_DFPRQX9 clk_r_REG176_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [27]), 
        .CP(clk), .RN(n9362), .Q(n8769) );
  HS65_LH_DFPRQX9 clk_r_REG125_S4 ( .D(\u_DataPath/pc4_to_idexreg_i [13]), 
        .CP(clk), .RN(n9362), .Q(n8803) );
  HS65_LH_DFPRQX9 clk_r_REG366_S3 ( .D(\u_DataPath/pc4_to_idexreg_i [1]), .CP(
        clk), .RN(n9362), .Q(n8808) );
  HS65_LH_DFPRQX9 clk_r_REG257_S3 ( .D(\u_DataPath/pc_4_i [12]), .CP(clk), 
        .RN(n9362), .Q(n9067) );
  HS65_LH_DFPRQX9 clk_r_REG169_S4 ( .D(\u_DataPath/pc_4_i [26]), .CP(clk), 
        .RN(n9362), .Q(n8976) );
  HS65_LH_DFPRQX9 clk_r_REG222_S3 ( .D(\u_DataPath/pc_4_i [19]), .CP(clk), 
        .RN(n9362), .Q(n8979) );
  HS65_LH_DFPRQX9 clk_r_REG235_S3 ( .D(\u_DataPath/pc_4_i [17]), .CP(clk), 
        .RN(n9362), .Q(n8994) );
  HS65_LH_DFPRQX9 clk_r_REG186_S4 ( .D(\u_DataPath/pc_4_i [30]), .CP(clk), 
        .RN(n9362), .Q(n8995) );
  HS65_LH_DFPRQX9 clk_r_REG614_S1 ( .D(n7923), .CP(clk), .RN(n9362), .Q(n9253)
         );
  HS65_LH_DFPRQX9 clk_r_REG539_S2 ( .D(n7920), .CP(clk), .RN(n9362), .Q(n9142)
         );
  HS65_LH_DFPRQX9 clk_r_REG618_S1 ( .D(iram_data[31]), .CP(clk), .RN(n9362), 
        .Q(n9333) );
  HS65_LH_DFPRQX9 clk_r_REG639_S1 ( .D(iram_data[7]), .CP(clk), .RN(n9362), 
        .Q(n9310) );
  HS65_LL_IVX18 U3679 ( .A(\u_DataPath/cw_towb_i [1]), .Z(n3030) );
  HS65_LH_IVX9 U4423 ( .A(n8968), .Z(n2947) );
  HS65_LH_DFPQNX4 clk_r_REG33_S1 ( .D(\u_DataPath/from_alu_data_out_i [8]), 
        .CP(clk), .QN(n3212) );
  HS65_LH_DFPQNX4 clk_r_REG109_S1 ( .D(\u_DataPath/from_alu_data_out_i [9]), 
        .CP(clk), .QN(n3079) );
  HS65_LH_DFPQNX4 clk_r_REG434_S1 ( .D(n8621), .CP(clk), .QN(n3016) );
  HS65_LL_DFPQNX4 clk_r_REG36_S1 ( .D(\u_DataPath/from_alu_data_out_i [11]), 
        .CP(clk), .QN(n3069) );
  HS65_LH_DFPQNX4 clk_r_REG90_S1 ( .D(\u_DataPath/from_alu_data_out_i [17]), 
        .CP(clk), .QN(n3024) );
  HS65_LH_DFPQNX4 clk_r_REG74_S1 ( .D(\u_DataPath/from_alu_data_out_i [13]), 
        .CP(clk), .QN(n3248) );
  HS65_LH_CBI4I1X5 U3841 ( .A(n8801), .B(n8893), .C(n9189), .D(n8432), .Z(
        \u_DataPath/dataOut_exe_i [3]) );
  HS65_LH_IVX18 U4322 ( .A(n9401), .Z(n2866) );
  HS65_LH_DFPQNX4 clk_r_REG15_S1 ( .D(\u_DataPath/from_alu_data_out_i [12]), 
        .CP(clk), .QN(n3259) );
  HS65_LL_DFPQNX4 clk_r_REG437_S1 ( .D(\u_DataPath/data_read_ex_2_i [3]), .CP(
        clk), .QN(n3309) );
  HS65_LH_DFPQNX4 clk_r_REG43_S1 ( .D(\u_DataPath/from_alu_data_out_i [31]), 
        .CP(clk), .QN(n3406) );
  HS65_LH_DFPQNX4 clk_r_REG21_S1 ( .D(\u_DataPath/from_alu_data_out_i [16]), 
        .CP(clk), .QN(n3093) );
  HS65_LH_DFPQNX4 clk_r_REG86_S1 ( .D(\u_DataPath/from_alu_data_out_i [22]), 
        .CP(clk), .QN(n3166) );
  HS65_LH_DFPQNX4 clk_r_REG18_S1 ( .D(\u_DataPath/from_alu_data_out_i [14]), 
        .CP(clk), .QN(n3088) );
  HS65_LH_DFPQNX4 clk_r_REG31_S1 ( .D(\u_DataPath/from_alu_data_out_i [30]), 
        .CP(clk), .QN(n3047) );
  HS65_LH_DFPQNX4 clk_r_REG94_S1 ( .D(\u_DataPath/from_alu_data_out_i [19]), 
        .CP(clk), .QN(n3185) );
  HS65_LH_DFPQNX4 clk_r_REG96_S1 ( .D(\u_DataPath/from_alu_data_out_i [20]), 
        .CP(clk), .QN(n3175) );
  HS65_LH_DFPQNX4 clk_r_REG293_S1 ( .D(n8579), .CP(clk), .QN(n2972) );
  HS65_LH_DFPQNX4 clk_r_REG40_S1 ( .D(\u_DataPath/from_alu_data_out_i [2]), 
        .CP(clk), .QN(n2934) );
  HS65_LH_DFPQNX4 clk_r_REG12_S1 ( .D(\u_DataPath/from_alu_data_out_i [7]), 
        .CP(clk), .QN(n3103) );
  HS65_LH_DFPQNX4 clk_r_REG64_S1 ( .D(\u_DataPath/from_alu_data_out_i [29]), 
        .CP(clk), .QN(n2968) );
  HS65_LH_DFPQNX4 clk_r_REG99_S1 ( .D(\u_DataPath/from_alu_data_out_i [23]), 
        .CP(clk), .QN(n3018) );
  HS65_LH_DFPQNX4 clk_r_REG103_S1 ( .D(\u_DataPath/u_memwbreg/N64 ), .CP(clk), 
        .QN(n7877) );
  HS65_LH_DFPQNX4 clk_r_REG105_S1 ( .D(\u_DataPath/from_alu_data_out_i [21]), 
        .CP(clk), .QN(n2956) );
  HS65_LH_DFPQNX4 clk_r_REG80_S1 ( .D(\u_DataPath/from_alu_data_out_i [24]), 
        .CP(clk), .QN(n3137) );
  HS65_LH_DFPQNX4 clk_r_REG7_S1 ( .D(\u_DataPath/from_alu_data_out_i [3]), 
        .CP(clk), .QN(n2970) );
  HS65_LH_DFPQNX4 clk_r_REG56_S1 ( .D(\u_DataPath/from_alu_data_out_i [5]), 
        .CP(clk), .QN(n3332) );
  HS65_LL_NAND2AX14 U3939 ( .A(n3289), .B(n2910), .Z(n5136) );
  HS65_LL_IVX18 U4300 ( .A(n3082), .Z(n3341) );
  HS65_LH_DFPQNX4 clk_r_REG25_S1 ( .D(\u_DataPath/from_alu_data_out_i [18]), 
        .CP(clk), .QN(n3084) );
  HS65_LH_DFPQNX4 clk_r_REG83_S1 ( .D(\u_DataPath/from_alu_data_out_i [25]), 
        .CP(clk), .QN(n3098) );
  HS65_LH_NAND3AX6 U3714 ( .A(n8507), .B(n9376), .C(n8508), .Z(n3245) );
  HS65_LH_IVX9 U3930 ( .A(n2845), .Z(n2855) );
  HS65_LL_DFPQNX4 clk_r_REG279_S1 ( .D(\u_DataPath/data_read_ex_2_i [26]), 
        .CP(clk), .QN(n3152) );
  HS65_LL_DFPQNX4 clk_r_REG341_S1 ( .D(\u_DataPath/data_read_ex_2_i [24]), 
        .CP(clk), .QN(n3143) );
  HS65_LL_DFPQNX4 clk_r_REG361_S1 ( .D(\u_DataPath/data_read_ex_1_i [5]), .CP(
        clk), .QN(n3335) );
  HS65_LL_DFPQNX4 clk_r_REG356_S2 ( .D(\u_DataPath/data_read_ex_2_i [28]), 
        .CP(clk), .QN(n3128) );
  HS65_LH_NAND2AX7 U4801 ( .A(n3058), .B(n2916), .Z(n4726) );
  HS65_LL_AOI21X2 U6685 ( .A(n4175), .B(n3237), .C(n3066), .Z(n3067) );
  HS65_LL_NAND2AX7 U3938 ( .A(n3068), .B(n3067), .Z(\sub_x_53/A[0] ) );
  HS65_LL_NOR2AX6 U6694 ( .A(n2913), .B(n3295), .Z(\sub_x_53/A[2] ) );
  HS65_LL_NOR2X6 U5629 ( .A(n3139), .B(n3138), .Z(\lte_x_59/B[24] ) );
  HS65_LL_IVX18 U3931 ( .A(n2845), .Z(n2856) );
  HS65_LL_IVX9 U4762 ( .A(n2855), .Z(n4587) );
  HS65_LH_IVX9 U3929 ( .A(n3432), .Z(n5004) );
  HS65_LH_NOR2X9 U3955 ( .A(n3474), .B(n5104), .Z(n3990) );
  HS65_LH_IVX9 U4755 ( .A(\lte_x_59/B[24] ), .Z(n4981) );
  HS65_LH_IVX9 U7378 ( .A(\lte_x_59/B[3] ), .Z(n5320) );
  HS65_LH_OAI12X3 U5426 ( .A(n3101), .B(n4795), .C(n3964), .Z(n4256) );
  HS65_LH_IVX9 U3607 ( .A(n4836), .Z(n4581) );
  HS65_LH_OAI12X3 U5416 ( .A(n2854), .B(n4795), .C(n3719), .Z(n4500) );
  HS65_LH_OAI12X3 U3713 ( .A(n4084), .B(n4081), .C(n4083), .Z(n4927) );
  HS65_LH_IVX9 U5614 ( .A(n7623), .Z(n7627) );
  HS65_LH_AOI21X2 U4124 ( .A(n3474), .B(n4587), .C(n3672), .Z(n3673) );
  HS65_LL_AND2X4 U3674 ( .A(n3356), .B(n3355), .Z(n3357) );
  HS65_LH_OAI12X3 U5525 ( .A(n4846), .B(n3558), .C(n3559), .Z(n5260) );
  HS65_LH_AOI21X2 U4105 ( .A(n2842), .B(n4587), .C(n3955), .Z(n3760) );
  HS65_LL_NOR2X6 U4183 ( .A(n2851), .B(n7627), .Z(n5342) );
  HS65_LH_AOI21X2 U7697 ( .A(n6035), .B(n5924), .C(n5923), .Z(n5925) );
  HS65_LH_IVX9 U4764 ( .A(n5201), .Z(n5131) );
  HS65_LL_NOR2X6 U4758 ( .A(n3818), .B(n4863), .Z(n5144) );
  HS65_LL_NOR2AX6 U5259 ( .A(n2867), .B(n3501), .Z(n5210) );
  HS65_LL_AOI21X2 U3893 ( .A(n4836), .B(n4491), .C(n4490), .Z(n4938) );
  HS65_LL_AOI21X2 U3962 ( .A(n4836), .B(n4840), .C(n4433), .Z(n4473) );
  HS65_LH_AOI21X2 U4039 ( .A(n5672), .B(n3598), .C(n3597), .Z(n3608) );
  HS65_LHS_XNOR2X3 U7745 ( .A(\u_DataPath/jaddr_i [22]), .B(n8966), .Z(n7104)
         );
  HS65_LL_XNOR2X4 U3786 ( .A(n8164), .B(n7086), .Z(n7080) );
  HS65_LHS_XNOR2X3 U7689 ( .A(n8165), .B(n2847), .Z(n7076) );
  HS65_LHS_XNOR2X3 U7663 ( .A(\u_DataPath/jaddr_i [18]), .B(n2847), .Z(n7085)
         );
  HS65_LH_DFPQNX9 clk_r_REG454_S1 ( .D(
        \u_DataPath/u_decode_unit/hdu_0/current_state [0]), .CP(clk), .QN(
        n7613) );
  HS65_LH_NOR2X6 U7651 ( .A(n6150), .B(n6139), .Z(n6634) );
  HS65_LH_NOR2X6 U3759 ( .A(n6150), .B(n6149), .Z(n6384) );
  HS65_LH_NOR2AX3 U6856 ( .A(n8729), .B(n3115), .Z(n2995) );
  HS65_LH_NOR2AX3 U3681 ( .A(n8736), .B(n2994), .Z(n8671) );
  HS65_LH_NOR2AX3 U3683 ( .A(n8737), .B(n2994), .Z(n8673) );
  HS65_LH_NOR2AX3 U3693 ( .A(n8727), .B(n2994), .Z(n8672) );
  HS65_LH_NOR2AX3 U3701 ( .A(n8874), .B(n2994), .Z(n3013) );
  HS65_LH_NOR2AX3 U3691 ( .A(\u_DataPath/dataOut_exe_i [11]), .B(n2986), .Z(
        n2993) );
  HS65_LH_NOR2AX3 U6775 ( .A(\u_DataPath/dataOut_exe_i [21]), .B(n3116), .Z(
        n3001) );
  HS65_LH_NOR2AX3 U6769 ( .A(\u_DataPath/dataOut_exe_i [22]), .B(n3116), .Z(
        n2989) );
  HS65_LH_NOR2AX3 U6770 ( .A(\u_DataPath/dataOut_exe_i [25]), .B(n3116), .Z(
        n2987) );
  HS65_LH_NOR2AX3 U6774 ( .A(\u_DataPath/dataOut_exe_i [24]), .B(n3116), .Z(
        n3004) );
  HS65_LH_NOR2AX3 U6777 ( .A(\u_DataPath/dataOut_exe_i [20]), .B(n3116), .Z(
        n3000) );
  HS65_LH_NOR2AX3 U6779 ( .A(\u_DataPath/dataOut_exe_i [30]), .B(n3116), .Z(
        n3002) );
  HS65_LH_AOI21X2 U6280 ( .A(n5284), .B(n5285), .C(n4302), .Z(n7839) );
  HS65_LL_NAND2X7 U3946 ( .A(n3204), .B(n3203), .Z(n5001) );
  HS65_LL_AOI12X2 U4319 ( .A(n6109), .B(n6111), .C(n5940), .Z(n6029) );
  HS65_LH_NOR2AX3 U6857 ( .A(n8749), .B(n3115), .Z(n2999) );
  HS65_LH_NOR2AX3 U6860 ( .A(n9241), .B(n3115), .Z(n2996) );
  HS65_LH_IVX9 U3434 ( .A(n8698), .Z(n9357) );
  HS65_LL_NOR2X6 U3437 ( .A(n6153), .B(n6149), .Z(n6317) );
  HS65_LL_AOI21X2 U3446 ( .A(\lte_x_59/B[18] ), .B(n4588), .C(n3954), .Z(n4258) );
  HS65_LL_NOR2X6 U3447 ( .A(n5152), .B(n4581), .Z(n4942) );
  HS65_LH_IVX18 U3448 ( .A(n5173), .Z(n5667) );
  HS65_LL_NAND2X7 U3465 ( .A(n4949), .B(n3426), .Z(n5173) );
  HS65_LL_OAI21X3 U3499 ( .A(n8427), .B(n9401), .C(n3135), .Z(n8554) );
  HS65_LL_IVX18 U3508 ( .A(n2893), .Z(n4351) );
  HS65_LL_NOR2X2 U3509 ( .A(n9401), .B(n8311), .Z(n8498) );
  HS65_LL_MUXI21X2 U3511 ( .D0(n2934), .D1(n2933), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8488) );
  HS65_LL_IVX18 U3512 ( .A(n9376), .Z(n4713) );
  HS65_LL_IVX18 U3516 ( .A(n3119), .Z(addr_to_iram[24]) );
  HS65_LH_IVX40 U3526 ( .A(n9357), .Z(addr_to_iram[11]) );
  HS65_LL_NAND2X7 U3538 ( .A(\u_DataPath/dataOut_exe_i [0]), .B(n3114), .Z(
        n8270) );
  HS65_LL_AOI12X9 U3540 ( .A(n5858), .B(n5860), .C(n5741), .Z(n5854) );
  HS65_LL_NOR2X6 U3547 ( .A(n6153), .B(n6132), .Z(n6624) );
  HS65_LL_OAI21X12 U3555 ( .A(n5743), .B(n5746), .C(n5745), .Z(n5860) );
  HS65_LL_AOI21X6 U3567 ( .A(n5285), .B(n3514), .C(n3513), .Z(n8479) );
  HS65_LL_NOR2AX3 U3570 ( .A(n5225), .B(n5224), .Z(n8458) );
  HS65_LL_NAND3X5 U3571 ( .A(n4416), .B(n2900), .C(n4415), .Z(n5166) );
  HS65_LL_AND3X4 U3572 ( .A(n4406), .B(n4405), .C(n4404), .Z(n2900) );
  HS65_LL_NAND2X7 U3575 ( .A(\u_DataPath/jaddr_i [23]), .B(n6131), .Z(n6132)
         );
  HS65_LL_AOI21X6 U3581 ( .A(n5285), .B(n4963), .C(n4962), .Z(n8475) );
  HS65_LH_NAND4ABX3 U3582 ( .A(n3845), .B(n3844), .C(n3843), .D(n3842), .Z(
        n3851) );
  HS65_LH_OAI21X3 U3584 ( .A(n5462), .B(n5461), .C(n5460), .Z(n5498) );
  HS65_LL_AOI21X2 U3585 ( .A(n5234), .B(n3610), .C(n3609), .Z(n3611) );
  HS65_LL_OAI12X3 U3587 ( .A(n2859), .B(n4324), .C(n4323), .Z(n4325) );
  HS65_LL_NOR4ABX2 U3591 ( .A(n4959), .B(n4958), .C(n4957), .D(n4956), .Z(
        n4960) );
  HS65_LL_NOR2AX3 U3593 ( .A(n5253), .B(n5252), .Z(n5268) );
  HS65_LH_AOI21X2 U3603 ( .A(n5667), .B(n5666), .C(n5665), .Z(n5668) );
  HS65_LH_AOI21X2 U3606 ( .A(n5667), .B(n4184), .C(n4183), .Z(n4202) );
  HS65_LH_OAI12X3 U3623 ( .A(n3246), .B(n3815), .C(n3950), .Z(n3951) );
  HS65_LH_NOR2AX3 U3624 ( .A(n5217), .B(n4936), .Z(n4961) );
  HS65_LH_NAND3X3 U3627 ( .A(n3608), .B(n2930), .C(n3607), .Z(n3609) );
  HS65_LH_AOI21X2 U3629 ( .A(n5618), .B(n4389), .C(n3600), .Z(n2930) );
  HS65_LL_OAI21X2 U3630 ( .A(n7634), .B(n9339), .C(n4126), .Z(n4139) );
  HS65_LH_AOI21X2 U3631 ( .A(n5667), .B(n5644), .C(n3784), .Z(n3785) );
  HS65_LL_NOR2AX3 U3633 ( .A(n5636), .B(n5635), .Z(n5637) );
  HS65_LL_AOI21X2 U3636 ( .A(n4480), .B(n4645), .C(n4102), .Z(n4103) );
  HS65_LH_AOI21X2 U3638 ( .A(n5667), .B(n5203), .C(n4434), .Z(n4444) );
  HS65_LH_AOI21X2 U3641 ( .A(n5618), .B(n5174), .C(n4436), .Z(n4443) );
  HS65_LL_AOI21X2 U3643 ( .A(n5629), .B(n3379), .C(n3378), .Z(n3380) );
  HS65_LL_AOI21X2 U3645 ( .A(n6123), .B(n5671), .C(n4168), .Z(n4169) );
  HS65_LL_AOI21X2 U3651 ( .A(n4259), .B(n4258), .C(n4581), .Z(n4261) );
  HS65_LL_NOR4ABX4 U3655 ( .A(n4125), .B(n4124), .C(n4123), .D(n4122), .Z(
        n4126) );
  HS65_LH_AOI21X2 U3659 ( .A(n3893), .B(n5294), .C(n5406), .Z(n5521) );
  HS65_LL_AOI21X2 U3663 ( .A(\sub_x_53/A[20] ), .B(n4544), .C(n3953), .Z(n4259) );
  HS65_LL_NOR2X6 U3664 ( .A(n4965), .B(n3416), .Z(n5285) );
  HS65_LH_AOI21X2 U3667 ( .A(\lte_x_59/B[22] ), .B(n4588), .C(n3779), .Z(n3780) );
  HS65_LH_NAND3X5 U3669 ( .A(n3837), .B(n3436), .C(n3435), .Z(n5170) );
  HS65_LH_AOI21X2 U3672 ( .A(n5667), .B(n5658), .C(n4166), .Z(n4167) );
  HS65_LL_CNIVX7 U3678 ( .A(n5249), .Z(n5672) );
  HS65_LL_AND2X4 U3682 ( .A(n4949), .B(n4508), .Z(n5661) );
  HS65_LL_NAND2AX14 U3689 ( .A(n2924), .B(n3492), .Z(n4879) );
  HS65_LL_OA12X9 U3694 ( .A(n4101), .B(n3358), .C(n3357), .Z(n3815) );
  HS65_LL_CNIVX7 U3708 ( .A(n5178), .Z(n5649) );
  HS65_LH_AOI21X2 U3712 ( .A(\lte_x_59/B[5] ), .B(n4544), .C(n3669), .Z(n3921)
         );
  HS65_LL_IVX9 U3722 ( .A(n3529), .Z(n5647) );
  HS65_LH_IVX27 U3737 ( .A(n3789), .Z(n4582) );
  HS65_LL_IVX9 U3741 ( .A(n4795), .Z(n3789) );
  HS65_LL_BFX9 U3751 ( .A(n2893), .Z(n5129) );
  HS65_LL_NAND2X21 U3753 ( .A(n3399), .B(n5136), .Z(n4795) );
  HS65_LL_IVX9 U3756 ( .A(n3430), .Z(n2872) );
  HS65_LH_IVX9 U3773 ( .A(n4147), .Z(n2865) );
  HS65_LL_NOR2X6 U3775 ( .A(n3417), .B(n3416), .Z(n3967) );
  HS65_LL_OAI12X6 U3776 ( .A(n3196), .B(n8531), .C(n3195), .Z(n5005) );
  HS65_LL_NAND2X7 U3777 ( .A(n3209), .B(n3208), .Z(n5021) );
  HS65_LH_NOR2X13 U3780 ( .A(n3306), .B(n3305), .Z(\lte_x_59/B[3] ) );
  HS65_LL_OAI12X6 U3781 ( .A(n3325), .B(n8498), .C(n3324), .Z(n4147) );
  HS65_LL_OAI21X3 U3798 ( .A(n8394), .B(n3340), .C(n3304), .Z(n3305) );
  HS65_LL_AOI21X2 U3803 ( .A(n3167), .B(n3270), .C(n2911), .Z(n3168) );
  HS65_LL_CNIVX7 U3807 ( .A(\u_DataPath/u_idexreg/N3 ), .Z(n7834) );
  HS65_LH_AOI21X2 U3813 ( .A(n2896), .B(n3134), .C(n3133), .Z(n3135) );
  HS65_LL_OAI12X6 U3819 ( .A(n3245), .B(n3244), .C(n3243), .Z(n5104) );
  HS65_LL_NAND4ABX3 U3820 ( .A(n8129), .B(n8892), .C(n8886), .D(n8126), .Z(
        \u_DataPath/u_idexreg/N3 ) );
  HS65_LL_MUXI21X5 U3825 ( .D0(n2970), .D1(n2969), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8394) );
  HS65_LL_MUXI21X2 U3831 ( .D0(n3332), .D1(n3331), .S0(n3404), .Z(n8391) );
  HS65_LH_OAI12X3 U3832 ( .A(n9190), .B(n8890), .C(n8317), .Z(
        \u_DataPath/dataOut_exe_i [26]) );
  HS65_LH_MUXI21X2 U3839 ( .D0(n8907), .D1(
        \u_DataPath/from_mem_data_out_i [10]), .S0(\u_DataPath/cw_towb_i [0]), 
        .Z(n8258) );
  HS65_LL_OAI12X3 U3843 ( .A(n8777), .B(n8114), .C(n8878), .Z(n8078) );
  HS65_LL_OAI21X2 U3845 ( .A(n8702), .B(n9012), .C(n8101), .Z(n8103) );
  HS65_LH_OAI12X3 U3849 ( .A(n9190), .B(n9072), .C(n8333), .Z(
        \u_DataPath/dataOut_exe_i [9]) );
  HS65_LL_OAI13X5 U3850 ( .A(n8904), .B(n9051), .C(n9081), .D(n8880), .Z(n8440) );
  HS65_LL_OAI12X3 U3852 ( .A(n9051), .B(n9103), .C(n8898), .Z(n8441) );
  HS65_LL_AOI21X6 U3863 ( .A(n9130), .B(n8750), .C(\u_DataPath/u_idexreg/N10 ), 
        .Z(n8071) );
  HS65_LL_OR3X9 U3866 ( .A(\u_DataPath/cw_exmem_i [5]), .B(
        \u_DataPath/cw_exmem_i [3]), .C(n9152), .Z(\u_DataPath/u_idexreg/N10 )
         );
  HS65_LH_IVX2 U3870 ( .A(n5056), .Z(n5057) );
  HS65_LH_OAI21X2 U3872 ( .A(n5123), .B(n5179), .C(n5137), .Z(n5138) );
  HS65_LH_NAND3X2 U3873 ( .A(n4971), .B(n4970), .C(n4969), .Z(n4972) );
  HS65_LH_NAND2X2 U3875 ( .A(n5144), .B(n5143), .Z(n5145) );
  HS65_LH_NAND2X2 U3876 ( .A(n5387), .B(n4143), .Z(n5550) );
  HS65_LH_IVX2 U3884 ( .A(n4997), .Z(n5345) );
  HS65_LH_NOR2X2 U3895 ( .A(n3285), .B(n4713), .Z(n3286) );
  HS65_LH_NAND2X2 U3904 ( .A(n4714), .B(n8557), .Z(n3154) );
  HS65_LH_IVX2 U3905 ( .A(n4750), .Z(n4752) );
  HS65_LH_IVX2 U3910 ( .A(n5550), .Z(n5551) );
  HS65_LH_IVX2 U3911 ( .A(n5313), .Z(n5107) );
  HS65_LH_IVX2 U3914 ( .A(n5035), .Z(n5549) );
  HS65_LH_IVX2 U3940 ( .A(n8528), .Z(n3202) );
  HS65_LH_NAND2X2 U3944 ( .A(n5320), .B(n5321), .Z(n5317) );
  HS65_LH_NAND2X2 U3956 ( .A(n4738), .B(n4737), .Z(n4747) );
  HS65_LH_NAND2X2 U3968 ( .A(n5323), .B(n5322), .Z(n5324) );
  HS65_LH_NAND2X2 U3976 ( .A(n5408), .B(n5378), .Z(n5412) );
  HS65_LH_NAND3X2 U3978 ( .A(n5322), .B(n5318), .C(n5317), .Z(n5332) );
  HS65_LH_IVX2 U3979 ( .A(n8559), .Z(n3146) );
  HS65_LH_AOI21X2 U3981 ( .A(n4351), .B(\sub_x_53/A[27] ), .C(n4350), .Z(n4353) );
  HS65_LH_IVX2 U3982 ( .A(n8516), .Z(n3251) );
  HS65_LH_NAND2X2 U3989 ( .A(n2849), .B(n4351), .Z(n3594) );
  HS65_LH_IVX2 U4002 ( .A(n5627), .Z(n5628) );
  HS65_LH_NAND2X2 U4011 ( .A(n4713), .B(n9030), .Z(n4655) );
  HS65_LH_NAND2X2 U4013 ( .A(n2842), .B(n2864), .Z(n3956) );
  HS65_LH_IVX2 U4023 ( .A(n5347), .Z(n5566) );
  HS65_LH_NAND2X2 U4036 ( .A(n5290), .B(n5362), .Z(n4702) );
  HS65_LH_OAI21X2 U4047 ( .A(n5523), .B(n5522), .C(n5521), .Z(n5524) );
  HS65_LH_IVX2 U4049 ( .A(n5333), .Z(n5309) );
  HS65_LL_IVX2 U4053 ( .A(n5209), .Z(n3619) );
  HS65_LH_NOR2X2 U4056 ( .A(n3657), .B(n3656), .Z(n4180) );
  HS65_LH_NAND2X2 U4069 ( .A(\lte_x_59/B[7] ), .B(n2845), .Z(n4154) );
  HS65_LH_OAI21X2 U4073 ( .A(n4524), .B(n4523), .C(n5229), .Z(n4525) );
  HS65_LH_NAND2X2 U4074 ( .A(n3327), .B(n9267), .Z(n3253) );
  HS65_LH_IVX2 U4080 ( .A(n4355), .Z(n4394) );
  HS65_LH_NOR2X2 U4084 ( .A(n5005), .B(\lte_x_59/B[18] ), .Z(n4250) );
  HS65_LH_IVX2 U4087 ( .A(n3875), .Z(n3878) );
  HS65_LH_NOR2X2 U4090 ( .A(n2854), .B(n2893), .Z(n3834) );
  HS65_LH_AOI21X2 U4103 ( .A(\sub_x_53/A[29] ), .B(n4544), .C(n3648), .Z(n3652) );
  HS65_LH_IVX2 U4114 ( .A(n3990), .Z(n4041) );
  HS65_LH_IVX2 U4115 ( .A(n5629), .Z(n3702) );
  HS65_LH_IVX2 U4119 ( .A(n3908), .Z(n3909) );
  HS65_LH_IVX2 U4129 ( .A(n4180), .Z(n4184) );
  HS65_LH_IVX2 U4135 ( .A(n4320), .Z(n3471) );
  HS65_LH_NAND2X2 U4140 ( .A(\lte_x_59/B[14] ), .B(n4588), .Z(n3985) );
  HS65_LHS_XNOR2X3 U4141 ( .A(\u_DataPath/jaddr_i [17]), .B(n8966), .Z(n7099)
         );
  HS65_LH_OAI21X2 U4152 ( .A(n4344), .B(n4343), .C(n4342), .Z(n4345) );
  HS65_LH_IVX2 U4157 ( .A(n3932), .Z(n3933) );
  HS65_LH_IVX2 U4160 ( .A(n4108), .Z(n4476) );
  HS65_LH_NAND2X2 U4171 ( .A(n3426), .B(n4840), .Z(n4841) );
  HS65_LH_AOI22X1 U4174 ( .A(n3474), .B(n4587), .C(n4551), .D(\lte_x_59/B[9] ), 
        .Z(n4128) );
  HS65_LH_OA12X4 U4178 ( .A(n4641), .B(n4637), .C(n4663), .Z(n3355) );
  HS65_LH_IVX2 U4189 ( .A(n5806), .Z(n5734) );
  HS65_LH_NOR2X2 U4192 ( .A(n2843), .B(n3756), .Z(n3672) );
  HS65_LH_NAND2X2 U4193 ( .A(n4824), .B(n3486), .Z(n4825) );
  HS65_LH_OAI21X2 U4198 ( .A(n4643), .B(n4642), .C(n4641), .Z(n4644) );
  HS65_LH_NAND2X2 U4202 ( .A(\lte_x_59/B[14] ), .B(n4544), .Z(n3832) );
  HS65_LH_NOR2X6 U4208 ( .A(n6353), .B(n6341), .Z(n6681) );
  HS65_LH_NAND2X2 U4231 ( .A(n4943), .B(n3426), .Z(n3981) );
  HS65_LH_IVX2 U4235 ( .A(n4389), .Z(n3539) );
  HS65_LH_OAI21X2 U4244 ( .A(n3762), .B(n4955), .C(n3761), .Z(n3797) );
  HS65_LH_NAND2X2 U4260 ( .A(n4926), .B(n4925), .Z(n4935) );
  HS65_LH_NAND2X2 U4261 ( .A(n4238), .B(n5194), .Z(n4240) );
  HS65_LH_OAI21X2 U4266 ( .A(n4391), .B(n4855), .C(n3581), .Z(n3592) );
  HS65_LH_NAND3X2 U4271 ( .A(n3426), .B(n4507), .C(n5615), .Z(n3654) );
  HS65_LH_AOI21X2 U4274 ( .A(n5780), .B(n5726), .C(n5725), .Z(n5759) );
  HS65_LH_OR2X4 U4281 ( .A(\sub_x_53/A[30] ), .B(n4966), .Z(n4211) );
  HS65_LH_NAND3X2 U4287 ( .A(n4347), .B(n4346), .C(n4345), .Z(n4348) );
  HS65_LH_NOR2X2 U4290 ( .A(n4052), .B(n3815), .Z(n4053) );
  HS65_LH_NAND2X4 U4292 ( .A(n3374), .B(n5271), .Z(n4420) );
  HS65_LH_NOR2X2 U4301 ( .A(n4134), .B(n5249), .Z(n5186) );
  HS65_LH_NAND2X2 U4307 ( .A(n7631), .B(n5638), .Z(n5639) );
  HS65_LH_OAI21X2 U4314 ( .A(n3874), .B(n5201), .C(n3873), .Z(n3882) );
  HS65_LL_NOR3X4 U4318 ( .A(n9150), .B(n9128), .C(n9051), .Z(n8439) );
  HS65_LH_NAND2X14 U4329 ( .A(n9251), .B(n8897), .Z(n8453) );
  HS65_LH_NAND2X2 U4331 ( .A(n3415), .B(n5321), .Z(n3818) );
  HS65_LH_XNOR2X4 U4346 ( .A(\u_DataPath/jaddr_i [17]), .B(n7086), .Z(n7088)
         );
  HS65_LH_AO22X4 U4353 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][2] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][2] ), .D(n7318), .Z(n6959) );
  HS65_LH_AO22X4 U4367 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][21] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][21] ), .D(
        n7586), .Z(n7588) );
  HS65_LH_AOI22X1 U4369 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][24] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][24] ), .Z(n7566)
         );
  HS65_LH_AO22X4 U4384 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][29] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][29] ), .Z(n7532)
         );
  HS65_LH_AOI22X1 U4388 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][28] ), .B(n7603), 
        .C(n6966), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][28] ), .Z(n7505)
         );
  HS65_LH_AOI22X1 U4390 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ), .B(n7604), 
        .C(n7334), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][20] ), .Z(n7484)
         );
  HS65_LH_AOI22X1 U4394 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][20] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ), .D(
        n2891), .Z(n7475) );
  HS65_LH_AOI22X1 U4396 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][27] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][27] ), .D(
        n2891), .Z(n7455) );
  HS65_LH_AO22X4 U4400 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][0] ), .B(n7429), 
        .C(n7310), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][0] ), .Z(n7431) );
  HS65_LH_AOI22X1 U4404 ( .A(n6745), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][3] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][3] ), .D(n7516), 
        .Z(n7394) );
  HS65_LH_AOI22X1 U4411 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][14] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][14] ), .D(
        n2889), .Z(n7373) );
  HS65_LH_AOI22X1 U4414 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][4] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ), .D(n2889), .Z(n7353) );
  HS65_LH_BFX4 U4415 ( .A(n6952), .Z(n7310) );
  HS65_LH_BFX4 U4426 ( .A(n6682), .Z(n7592) );
  HS65_LH_NOR2X5 U4429 ( .A(n6148), .B(n6152), .Z(n2884) );
  HS65_LH_BFX4 U4453 ( .A(n6624), .Z(n6600) );
  HS65_LH_AOI22X1 U4473 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][2] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][2] ), .D(
        n6171), .Z(n6564) );
  HS65_LH_AO22X4 U4482 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][25] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][25] ), .D(
        n6629), .Z(n7147) );
  HS65_LH_AO22X4 U4485 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][9] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ), .D(n7291), .Z(n7138) );
  HS65_LH_AO22X4 U4486 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][28] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][28] ), .D(
        n7267), .Z(n6907) );
  HS65_LH_AO22X4 U4488 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][17] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][17] ), .D(
        n7267), .Z(n6887) );
  HS65_LH_AOI22X1 U4506 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][31] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][31] ), .D(
        n7272), .Z(n6873) );
  HS65_LH_AO22X4 U4507 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][18] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][18] ), .D(
        n7274), .Z(n6655) );
  HS65_LH_AO22X4 U4516 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][20] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][20] ), .D(
        n7276), .Z(n6851) );
  HS65_LH_AO22X4 U4526 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][5] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][5] ), .D(
        n7282), .Z(n6940) );
  HS65_LH_AO22X4 U4528 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][29] ), .D(
        n7282), .Z(n7290) );
  HS65_LH_AOI22X1 U4540 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][8] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ), .Z(n6776)
         );
  HS65_LH_AOI22X1 U4544 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][11] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][11] ), .D(
        n7285), .Z(n6254) );
  HS65_LH_AOI22X1 U4547 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][31] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][31] ), .Z(n6686)
         );
  HS65_LH_AOI22X1 U4548 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][25] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][25] ), .Z(n7049)
         );
  HS65_LH_AO22X4 U4549 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][6] ), .B(n7429), 
        .C(n7310), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][6] ), .Z(n7245) );
  HS65_LH_AOI22X1 U4554 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][21] ), .B(n6377), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][21] ), .D(
        n7171), .Z(n6193) );
  HS65_LH_AOI22X1 U4556 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][21] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ), .D(
        n6624), .Z(n6192) );
  HS65_LH_AOI22X1 U4557 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][16] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][16] ), .D(
        n6625), .Z(n6169) );
  HS65_LH_AO22X4 U4561 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][23] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][23] ), .D(
        n7318), .Z(n7229) );
  HS65_LH_AO22X4 U4585 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][1] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][1] ), .Z(n6838)
         );
  HS65_LH_AO22X4 U4596 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][27] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][27] ), .D(
        n6637), .Z(n6215) );
  HS65_LH_AOI22X1 U4600 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][19] ), .B(n7525), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ), .Z(n6755)
         );
  HS65_LH_AOI22X1 U4601 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][7] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][7] ), .Z(n6728)
         );
  HS65_LH_AO22X4 U4603 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][22] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][22] ), .D(
        n7292), .Z(n6279) );
  HS65_LH_AO22X4 U4614 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][24] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][24] ), .D(
        n7292), .Z(n6299) );
  HS65_LH_AO22X4 U4616 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][5] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][5] ), .Z(n6709)
         );
  HS65_LH_AOI22X1 U4619 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][5] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][5] ), .D(
        n6670), .Z(n6702) );
  HS65_LH_AO22X4 U4620 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][13] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][13] ), .D(
        n7292), .Z(n7178) );
  HS65_LH_AOI22X1 U4629 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][13] ), .B(n7165), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][13] ), .D(
        n6624), .Z(n7169) );
  HS65_LH_AOI22X1 U4634 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][14] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][14] ), .D(
        n6625), .Z(n6311) );
  HS65_LH_AO22X4 U4637 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][19] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][19] ), .D(
        n7267), .Z(n6515) );
  HS65_LH_AO22X4 U4643 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][7] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ), .D(n7267), .Z(n6435) );
  HS65_LH_AO22X4 U4659 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][12] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][12] ), .D(
        n7267), .Z(n6535) );
  HS65_LH_AO22X4 U4665 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][6] ), .B(n7275), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][6] ), .D(
        n7274), .Z(n6480) );
  HS65_LH_AO22X4 U4674 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ), .B(n6626), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[30][3] ), .D(
        n7274), .Z(n6580) );
  HS65_LH_AO22X4 U4678 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][26] ), .D(
        n7282), .Z(n6506) );
  HS65_LH_AO22X4 U4685 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][8] ), .B(n7283), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[20][8] ), .D(
        n7282), .Z(n6466) );
  HS65_LH_AOI22X1 U4691 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][1] ), .D(
        n7171), .Z(n6605) );
  HS65_LH_AOI22X1 U4697 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][11] ), .B(n7603), 
        .C(n7333), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ), .Z(n7069)
         );
  HS65_LH_NOR2AX3 U4707 ( .A(n3069), .B(\u_DataPath/cw_towb_i [0]), .Z(n3070)
         );
  HS65_LH_AO22X4 U4708 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][13] ), .B(n7578), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][13] ), .Z(n6977)
         );
  HS65_LH_AO22X4 U4712 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][22] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][22] ), .Z(n6996)
         );
  HS65_LH_AO22X4 U4713 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][4] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][4] ), .D(n7267), .Z(n6620) );
  HS65_LH_IVX2 U4715 ( .A(n3050), .Z(n3034) );
  HS65_LH_IVX2 U4723 ( .A(n4579), .Z(n4615) );
  HS65_LH_NOR2X2 U4742 ( .A(n4939), .B(n3979), .Z(n3989) );
  HS65_LH_IVX2 U4744 ( .A(n3515), .Z(n5293) );
  HS65_LH_IVX2 U4771 ( .A(n3698), .Z(n3699) );
  HS65_LH_NOR2X3 U4780 ( .A(\sub_x_53/A[2] ), .B(n3415), .Z(n4575) );
  HS65_LH_AOI21X2 U4786 ( .A(n4949), .B(n4948), .C(n4947), .Z(n4958) );
  HS65_LH_OAI21X2 U4792 ( .A(n5760), .B(n5878), .C(n5759), .Z(n5791) );
  HS65_LH_IVX2 U4799 ( .A(n5795), .Z(n5796) );
  HS65_LH_OR2X4 U4808 ( .A(n9342), .B(n9216), .Z(n5902) );
  HS65_LH_IVX2 U4814 ( .A(n5907), .Z(n5740) );
  HS65_LH_NAND2X2 U4817 ( .A(n9185), .B(n9230), .Z(n5789) );
  HS65_LH_NOR2X2 U4831 ( .A(n7645), .B(n7680), .Z(n7646) );
  HS65_LH_NOR2X2 U4833 ( .A(n9173), .B(n9231), .Z(n5874) );
  HS65_LH_NAND2X2 U4837 ( .A(n4050), .B(n3267), .Z(n4056) );
  HS65_LH_NAND2X2 U4843 ( .A(n5217), .B(n4885), .Z(n4900) );
  HS65_LH_IVX2 U4860 ( .A(n8262), .Z(n2966) );
  HS65_LH_NOR3X1 U4863 ( .A(\u_DataPath/dataOut_exe_i [1]), .B(n8360), .C(
        n8270), .Z(n7344) );
  HS65_LH_NAND2X2 U4872 ( .A(n5867), .B(n5866), .Z(n5869) );
  HS65_LH_OAI22X1 U4874 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [26]), .C(
        n8316), .D(n3409), .Z(n3151) );
  HS65_LH_NAND2X2 U4878 ( .A(n4713), .B(n9342), .Z(n4191) );
  HS65_LH_NAND2X2 U4886 ( .A(n9368), .B(n9008), .Z(n8435) );
  HS65_LH_NAND2X2 U4888 ( .A(n8687), .B(n8686), .Z(n7668) );
  HS65_LH_IVX2 U4906 ( .A(n8255), .Z(n3260) );
  HS65_LH_IVX2 U4909 ( .A(\u_DataPath/dataOut_exe_i [17]), .Z(n3201) );
  HS65_LH_AOI22X1 U4917 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][15] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][15] ), .Z(n7193)
         );
  HS65_LH_AO22X4 U4925 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][10] ), .B(n7523), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][10] ), .Z(n7214)
         );
  HS65_LH_AO22X4 U4927 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][0] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][0] ), .D(n7291), .Z(n6430) );
  HS65_LH_AOI22X1 U4928 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][10] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][10] ), .D(
        n7294), .Z(n6407) );
  HS65_LH_AOI22X1 U4936 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][15] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][15] ), .D(
        n6942), .Z(n6386) );
  HS65_LH_AOI22X1 U4938 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][15] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][15] ), .D(
        n7264), .Z(n6369) );
  HS65_LH_MUXI21X2 U4942 ( .D0(n2968), .D1(n9384), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8426) );
  HS65_LH_AOI21X2 U4948 ( .A(n3404), .B(n9386), .C(n3070), .Z(n8345) );
  HS65_LH_NAND2X2 U4956 ( .A(n9068), .B(n7773), .Z(n7690) );
  HS65_LH_OAI21X2 U4967 ( .A(n4255), .B(n4254), .C(n4516), .Z(n4265) );
  HS65_LH_IVX2 U4976 ( .A(n8056), .Z(n7698) );
  HS65_LH_IVX2 U4977 ( .A(n4538), .Z(n4574) );
  HS65_LL_OA12X4 U4982 ( .A(n7634), .B(n2844), .C(n4169), .Z(n4170) );
  HS65_LH_AOI22X1 U4986 ( .A(n8868), .B(n9029), .C(n9369), .D(n8939), .Z(n7845) );
  HS65_LH_NAND2X2 U4999 ( .A(n5777), .B(n5977), .Z(n5785) );
  HS65_LH_AOI21X2 U5004 ( .A(n5802), .B(n5868), .C(n5801), .Z(n5803) );
  HS65_LH_OAI21X2 U5005 ( .A(n6049), .B(n6045), .C(n6047), .Z(n6051) );
  HS65_LH_IVX2 U5013 ( .A(n5980), .Z(n5983) );
  HS65_LH_IVX2 U5015 ( .A(n6000), .Z(n6001) );
  HS65_LH_NAND2X2 U5016 ( .A(n7707), .B(n4003), .Z(n4287) );
  HS65_LH_MUXI21X5 U5017 ( .D0(n3137), .D1(n9389), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8550) );
  HS65_LH_NAND2X2 U5032 ( .A(n3201), .B(n3407), .Z(n3198) );
  HS65_LH_AOI22X1 U5040 ( .A(n4951), .B(n4578), .C(n5667), .D(n5239), .Z(n4010) );
  HS65_LH_NOR2X2 U5046 ( .A(n8845), .B(n3341), .Z(n3169) );
  HS65_LH_OAI22X1 U5047 ( .A(n3264), .B(\u_DataPath/dataOut_exe_i [25]), .C(
        n8427), .D(n3409), .Z(n3099) );
  HS65_LH_NOR2AX3 U5050 ( .A(n8726), .B(n2994), .Z(n8675) );
  HS65_LH_NOR2AX3 U5057 ( .A(n8742), .B(n2994), .Z(n8674) );
  HS65_LH_NOR2AX3 U5092 ( .A(\u_DataPath/dataOut_exe_i [8]), .B(n2986), .Z(
        n3006) );
  HS65_LH_NOR2AX3 U5096 ( .A(\u_DataPath/dataOut_exe_i [23]), .B(n3116), .Z(
        n3003) );
  HS65_LH_IVX2 U5104 ( .A(n9112), .Z(n2984) );
  HS65_LH_AO22X4 U5115 ( .A(n9262), .B(n9188), .C(n9133), .D(n8982), .Z(
        \u_DataPath/jump_address_i [19]) );
  HS65_LH_AO22X4 U5122 ( .A(n9104), .B(n9188), .C(n9133), .D(n8951), .Z(
        \u_DataPath/jump_address_i [10]) );
  HS65_LH_IVX2 U5129 ( .A(n7668), .Z(n7743) );
  HS65_LH_NAND2X2 U5132 ( .A(n2985), .B(n3109), .Z(n8425) );
  HS65_LH_NAND2X2 U5133 ( .A(n3412), .B(n2866), .Z(n8491) );
  HS65_LH_NAND2X2 U5134 ( .A(n4208), .B(n7869), .Z(n8569) );
  HS65_LH_NAND2X2 U5136 ( .A(n3278), .B(n7869), .Z(n8521) );
  HS65_LL_NAND3X2 U5141 ( .A(n4511), .B(n4510), .C(n4509), .Z(n5248) );
  HS65_LH_OA12X4 U5143 ( .A(n4829), .B(n9402), .C(n4827), .Z(n2926) );
  HS65_LH_NOR4ABX2 U5144 ( .A(n6826), .B(n6825), .C(n6824), .D(n6823), .Z(
        n8175) );
  HS65_LH_NOR4ABX2 U5151 ( .A(n6718), .B(n6717), .C(n6716), .D(n6715), .Z(
        n8171) );
  HS65_LH_AOI31X2 U5152 ( .A(n4608), .B(n4607), .C(n4606), .D(n5152), .Z(n4653) );
  HS65_LH_BFX4 U5153 ( .A(n7306), .Z(n7917) );
  HS65_LH_NOR2X2 U5154 ( .A(n7641), .B(n7640), .Z(n8135) );
  HS65_LH_NOR2X2 U5155 ( .A(n5696), .B(n5695), .Z(n7118) );
  HS65_LH_OAI21X2 U5160 ( .A(n5967), .B(n6007), .C(n5966), .Z(n6059) );
  HS65_LH_NAND2X2 U5162 ( .A(n6076), .B(n6031), .Z(n6032) );
  HS65_LH_NOR2X2 U5164 ( .A(n7758), .B(n7757), .Z(n7663) );
  HS65_LH_NAND2X2 U5176 ( .A(n8708), .B(n7764), .Z(n7765) );
  HS65_LH_NAND2X2 U5181 ( .A(n6054), .B(n6053), .Z(n6056) );
  HS65_LH_NOR2X2 U5187 ( .A(n7793), .B(n7792), .Z(n7731) );
  HS65_LH_NAND2X2 U5196 ( .A(n5949), .B(n5948), .Z(n5951) );
  HS65_LH_IVX2 U5200 ( .A(n6034), .Z(n6095) );
  HS65_LH_NOR2X2 U5212 ( .A(n7697), .B(n7694), .Z(n8040) );
  HS65_LH_NOR2X2 U5221 ( .A(n4475), .B(n4474), .Z(n4487) );
  HS65_LH_AOI21X2 U5227 ( .A(n5667), .B(n4872), .C(n4871), .Z(n4912) );
  HS65_LH_NOR2X2 U5228 ( .A(\u_DataPath/dataOut_exe_i [10]), .B(n3264), .Z(
        n3240) );
  HS65_LH_OAI211X1 U5230 ( .A(n8302), .B(n8575), .C(n7346), .D(n7345), .Z(
        n8298) );
  HS65_LH_NAND3X2 U5232 ( .A(n9113), .B(n2984), .C(n7639), .Z(n3109) );
  HS65_LH_NAND2AX4 U5241 ( .A(n9031), .B(n7733), .Z(n8144) );
  HS65_LH_NAND2X4 U5246 ( .A(n7851), .B(n9061), .Z(
        \u_DataPath/dataOut_exe_i [16]) );
  HS65_LH_AO22X4 U5247 ( .A(n9254), .B(n8768), .C(n9132), .D(n9009), .Z(
        \u_DataPath/pc4_to_idexreg_i [4]) );
  HS65_LH_AO22X4 U5251 ( .A(n8786), .B(n9139), .C(n9333), .D(n9154), .Z(
        opcode_i[5]) );
  HS65_LH_NOR4ABX2 U5252 ( .A(n7203), .B(n7202), .C(n7201), .D(n7200), .Z(
        n8305) );
  HS65_LH_AO22X4 U5253 ( .A(n9254), .B(n8769), .C(n9240), .D(n9070), .Z(
        \u_DataPath/pc4_to_idexreg_i [27]) );
  HS65_LH_AO22X4 U5256 ( .A(n8780), .B(n9252), .C(n9307), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [4]) );
  HS65_LH_AO22X4 U5262 ( .A(n9254), .B(n8804), .C(n9240), .D(n8974), .Z(
        \u_DataPath/pc4_to_idexreg_i [10]) );
  HS65_LH_AO22X4 U5265 ( .A(n9254), .B(n8827), .C(n9240), .D(n9108), .Z(
        \u_DataPath/pc4_to_idexreg_i [31]) );
  HS65_LHS_XOR2X3 U5271 ( .A(n5946), .B(n5945), .Z(
        \u_DataPath/u_execute/resAdd1_i [31]) );
  HS65_LH_NAND2X2 U5275 ( .A(\u_DataPath/immediate_ext_dec_i [0]), .B(
        \u_DataPath/immediate_ext_dec_i [1]), .Z(n8092) );
  HS65_LHS_XNOR2X3 U5278 ( .A(n2782), .B(n7663), .Z(\u_DataPath/pc_4_i [19])
         );
  HS65_LHS_XNOR2X3 U5286 ( .A(n3124), .B(n7679), .Z(\u_DataPath/pc_4_i [17])
         );
  HS65_LHS_XNOR2X3 U5292 ( .A(n6092), .B(n6091), .Z(
        \u_DataPath/u_execute/resAdd1_i [7]) );
  HS65_LL_NOR2AX6 U5302 ( .A(n4369), .B(n4368), .Z(n8469) );
  HS65_LHS_XOR2X3 U5303 ( .A(n7783), .B(n7782), .Z(
        \u_DataPath/u_execute/link_value_i [9]) );
  HS65_LHS_XNOR2X3 U5304 ( .A(n2825), .B(n7704), .Z(\u_DataPath/pc_4_i [27])
         );
  HS65_LH_IVX2 U5307 ( .A(Data_out_fromRAM[20]), .Z(n8410) );
  HS65_LH_IVX2 U5316 ( .A(Data_out_fromRAM[21]), .Z(n8365) );
  HS65_LH_IVX2 U5318 ( .A(n7740), .Z(n8095) );
  HS65_LH_NOR2X2 U5323 ( .A(n9175), .B(n9227), .Z(n6085) );
  HS65_LH_IVX2 U5325 ( .A(n5882), .Z(n5883) );
  HS65_LH_NOR2X2 U5338 ( .A(n9145), .B(n9224), .Z(n5753) );
  HS65_LH_IVX2 U5340 ( .A(n5957), .Z(n5958) );
  HS65_LH_NOR2X2 U5342 ( .A(n9033), .B(n9215), .Z(n5894) );
  HS65_LH_IVX2 U5348 ( .A(n6097), .Z(n6098) );
  HS65_LH_NOR2X2 U5353 ( .A(n9179), .B(n9225), .Z(n6090) );
  HS65_LH_IVX2 U5363 ( .A(n5887), .Z(n5831) );
  HS65_LH_NOR2X2 U5365 ( .A(n8913), .B(n9219), .Z(n6041) );
  HS65_LH_IVX2 U5366 ( .A(n5839), .Z(n5890) );
  HS65_LH_OR2X4 U5370 ( .A(n6148), .B(n6151), .Z(n9335) );
  HS65_LH_OR2X4 U5372 ( .A(n9002), .B(n8751), .Z(n9336) );
  HS65_LH_OR2X4 U5391 ( .A(n9344), .B(n9345), .Z(n9337) );
  HS65_LH_NOR2X2 U5393 ( .A(n9267), .B(n9228), .Z(n5987) );
  HS65_LH_IVX2 U5403 ( .A(n5786), .Z(n5787) );
  HS65_LH_IVX2 U5404 ( .A(n5960), .Z(n6057) );
  HS65_LH_NAND2X2 U5411 ( .A(n9181), .B(n9226), .Z(n6058) );
  HS65_LH_IVX2 U5418 ( .A(n5863), .Z(n5764) );
  HS65_LH_NOR2X2 U5422 ( .A(n9039), .B(n9116), .Z(n5899) );
  HS65_LH_IVX2 U5428 ( .A(n6102), .Z(n6050) );
  HS65_LH_IVX2 U5438 ( .A(n5836), .Z(n5837) );
  HS65_LH_NOR2X2 U5443 ( .A(n9177), .B(n9229), .Z(n5879) );
  HS65_LH_IVX2 U5446 ( .A(n6078), .Z(n6031) );
  HS65_LH_NAND2X2 U5450 ( .A(n9171), .B(n9214), .Z(n5871) );
  HS65_LH_IVX2 U5452 ( .A(n6070), .Z(n5984) );
  HS65_LH_NOR2X2 U5454 ( .A(n9171), .B(n9214), .Z(n5778) );
  HS65_LH_IVX2 U5460 ( .A(n5979), .Z(n6069) );
  HS65_LH_NAND2X2 U5463 ( .A(n8913), .B(n9219), .Z(n5891) );
  HS65_LH_IVX2 U5466 ( .A(n6094), .Z(n6042) );
  HS65_LH_IVX2 U5467 ( .A(n5285), .Z(n4829) );
  HS65_LH_NOR2X2 U5469 ( .A(n9183), .B(n9232), .Z(n5775) );
  HS65_LH_IVX2 U5472 ( .A(n5976), .Z(n5977) );
  HS65_LH_IVX2 U5477 ( .A(n5789), .Z(n5790) );
  HS65_LH_NOR2X2 U5485 ( .A(n9185), .B(n9230), .Z(n5772) );
  HS65_LH_IVX2 U5494 ( .A(n5990), .Z(n6005) );
  HS65_LH_NOR2X2 U5497 ( .A(n9037), .B(n9212), .Z(n5846) );
  HS65_LH_IVX2 U5498 ( .A(n6045), .Z(n6046) );
  HS65_LH_NOR2X2 U5499 ( .A(n9173), .B(n9231), .Z(n6073) );
  HS65_LH_IVX2 U5501 ( .A(n5874), .Z(n5875) );
  HS65_LH_OA12X4 U5502 ( .A(n3899), .B(n3815), .C(n3898), .Z(n9338) );
  HS65_LHS_XNOR2X3 U5509 ( .A(n4111), .B(n4110), .Z(n9339) );
  HS65_LH_IVX9 U5510 ( .A(n8876), .Z(n9340) );
  HS65_LH_IVX9 U5514 ( .A(n9340), .Z(n9341) );
  HS65_LH_IVX9 U5516 ( .A(n9340), .Z(n9342) );
  HS65_LH_IVX9 U5520 ( .A(n9340), .Z(n9343) );
  HS65_LH_NOR2X2 U5521 ( .A(n9336), .B(n9337), .Z(\u_DataPath/cw_to_ex_i [15])
         );
  HS65_LH_CNIVX3 U5523 ( .A(n9347), .Z(n9344) );
  HS65_LH_CNIVX3 U5527 ( .A(n9146), .Z(n9345) );
  HS65_LH_IVX2 U5529 ( .A(n3582), .Z(n9346) );
  HS65_LL_NOR2X6 U5566 ( .A(n5491), .B(n3423), .Z(n3582) );
  HS65_LH_IVX9 U5570 ( .A(n3582), .Z(n4548) );
  HS65_LH_AOI21X6 U5581 ( .A(n5643), .B(n4861), .C(n2902), .Z(n4862) );
  HS65_LL_BFX9 U5584 ( .A(n5179), .Z(n9348) );
  HS65_LH_AOI12X3 U5591 ( .A(n9349), .B(n5005), .C(n5649), .Z(n4269) );
  HS65_LH_NAND3X5 U5610 ( .A(n4990), .B(n5115), .C(n4989), .Z(n4991) );
  HS65_LL_IVX2 U5617 ( .A(n5082), .Z(n5529) );
  HS65_LH_NOR2X2 U5625 ( .A(n8824), .B(n3403), .Z(n3086) );
  HS65_LH_OAI21X2 U5637 ( .A(n4905), .B(n3815), .C(n5397), .Z(n4906) );
  HS65_LH_IVX7 U5658 ( .A(n9330), .Z(n9354) );
  HS65_LH_IVX7 U5660 ( .A(n9330), .Z(n9355) );
  HS65_LH_IVX7 U5664 ( .A(n9330), .Z(n9356) );
  HS65_LHS_XOR2X3 U5678 ( .A(addr_to_iram[29]), .B(n7786), .Z(
        \u_DataPath/pc_4_i [31]) );
  HS65_LH_IVX44 U5688 ( .A(n2780), .Z(addr_to_iram[29]) );
  HS65_LH_IVX44 U5691 ( .A(n3124), .Z(addr_to_iram[15]) );
  HS65_LH_IVX2 U5704 ( .A(n8677), .Z(n9359) );
  HS65_LH_IVX4 U5713 ( .A(n9359), .Z(n9360) );
  HS65_LH_IVX7 U5715 ( .A(n9359), .Z(n9361) );
  HS65_LH_IVX4 U5731 ( .A(n9359), .Z(n9362) );
  HS65_LH_IVX9 U5760 ( .A(n9135), .Z(n9364) );
  HS65_LH_IVX9 U5778 ( .A(n9364), .Z(n9365) );
  HS65_LH_IVX9 U5811 ( .A(n9364), .Z(n9366) );
  HS65_LH_IVX9 U5815 ( .A(n9135), .Z(n9367) );
  HS65_LH_IVX9 U5816 ( .A(n9367), .Z(n9368) );
  HS65_LH_IVX9 U5826 ( .A(n9367), .Z(n9369) );
  HS65_LH_AOI21X2 U5836 ( .A(n9007), .B(n9347), .C(n8082), .Z(n8088) );
  HS65_LL_OR2X18 U5854 ( .A(n3401), .B(n5136), .Z(n2893) );
  HS65_LH_OAI21X2 U5866 ( .A(n3427), .B(n5620), .C(n3767), .Z(n3795) );
  HS65_LH_OAI21X3 U5874 ( .A(n5173), .B(n5620), .C(n3986), .Z(n3987) );
  HS65_LL_NAND3X5 U5887 ( .A(n2931), .B(n4048), .C(n4047), .Z(n4302) );
  HS65_LH_OAI21X2 U5890 ( .A(n2848), .B(n3756), .C(n4154), .Z(n4155) );
  HS65_LH_NAND2X7 U5894 ( .A(n5643), .B(n4046), .Z(n4047) );
  HS65_LH_IVX9 U5895 ( .A(n5088), .Z(n3415) );
  HS65_LL_NAND4ABX6 U5914 ( .A(n5601), .B(n5600), .C(n8460), .D(n5599), .Z(
        n5678) );
  HS65_LL_AOI12X2 U5930 ( .A(n5415), .B(n5414), .C(n5413), .Z(n5462) );
  HS65_LH_AOI21X6 U5939 ( .A(n5459), .B(n5458), .C(n5457), .Z(n5460) );
  HS65_LH_NOR2X6 U5940 ( .A(\sub_x_53/A[27] ), .B(n3385), .Z(n3629) );
  HS65_LL_IVX2 U5942 ( .A(n4976), .Z(n3385) );
  HS65_LL_NAND2X2 U5957 ( .A(n4714), .B(n8546), .Z(n3171) );
  HS65_LL_NOR3AX9 U5959 ( .A(n4456), .B(n4455), .C(n4454), .Z(n5681) );
  HS65_LL_AOI21X2 U5963 ( .A(n4295), .B(n5211), .C(n4294), .Z(n4299) );
  HS65_LL_NAND2AX14 U5967 ( .A(n3381), .B(n3380), .Z(n5195) );
  HS65_LL_CNIVX3 U5970 ( .A(n5714), .Z(n4788) );
  HS65_LL_NOR3X7 U5978 ( .A(n4787), .B(n4786), .C(n4785), .Z(n5714) );
  HS65_LL_NAND3X3 U5982 ( .A(n2919), .B(n3202), .C(n8529), .Z(n3203) );
  HS65_LL_OAI12X6 U5986 ( .A(n3501), .B(n4426), .C(n3500), .Z(n5211) );
  HS65_LL_NOR2X2 U6012 ( .A(\sub_x_53/A[27] ), .B(n4976), .Z(n3682) );
  HS65_LL_OAI21X2 U6015 ( .A(n4736), .B(n4735), .C(n4734), .Z(n4783) );
  HS65_LL_BFX4 U6018 ( .A(n6618), .Z(n9370) );
  HS65_LH_BFX9 U6024 ( .A(n6618), .Z(n9371) );
  HS65_LH_BFX2 U6030 ( .A(n6618), .Z(n9372) );
  HS65_LL_NOR2X2 U6031 ( .A(n6148), .B(n6149), .Z(n6618) );
  HS65_LL_AOI22X3 U6034 ( .A(\lte_x_59/B[1] ), .B(n4588), .C(n4587), .D(
        \sub_x_53/A[0] ), .Z(n4117) );
  HS65_LH_BFX9 U6039 ( .A(n7312), .Z(n9373) );
  HS65_LH_NOR2X2 U6053 ( .A(n6353), .B(n6331), .Z(n7312) );
  HS65_LH_NOR2X2 U6060 ( .A(n5530), .B(n3515), .Z(n5416) );
  HS65_LH_NAND2X7 U6070 ( .A(n3420), .B(n4512), .Z(n5178) );
  HS65_LH_AOI12X3 U6087 ( .A(n5207), .B(n5658), .C(n4271), .Z(n4272) );
  HS65_LH_AOI21X2 U6094 ( .A(n4051), .B(n4918), .C(n5476), .Z(n4054) );
  HS65_LL_NAND2AX7 U6097 ( .A(n3364), .B(n3363), .Z(n4918) );
  HS65_LL_AOI21X2 U6113 ( .A(n5195), .B(n4335), .C(n4334), .Z(n4336) );
  HS65_LL_NOR2AX6 U6115 ( .A(n3387), .B(n3386), .Z(n4332) );
  HS65_LL_OAI21X2 U6116 ( .A(n3749), .B(n3629), .C(n5443), .Z(n3386) );
  HS65_LL_NOR2X6 U6118 ( .A(\lte_x_59/B[15] ), .B(n4677), .Z(n3891) );
  HS65_LH_IVX9 U6121 ( .A(n3891), .Z(n3892) );
  HS65_LH_NOR2X6 U6122 ( .A(n3891), .B(n4913), .Z(n3368) );
  HS65_LH_OAI12X3 U6126 ( .A(n5435), .B(n3698), .C(n3700), .Z(n3378) );
  HS65_LH_OAI21X2 U6131 ( .A(n4671), .B(n4583), .C(n4060), .Z(n4078) );
  HS65_LH_OAI22X1 U6132 ( .A(n2848), .B(n4583), .C(n3756), .D(n5041), .Z(n4130) );
  HS65_LH_OA12X4 U6134 ( .A(n5652), .B(n4583), .C(n3550), .Z(n2899) );
  HS65_LH_OAI22X1 U6135 ( .A(n5652), .B(n4583), .C(n3756), .D(n2860), .Z(n3666) );
  HS65_LL_NOR2X2 U6136 ( .A(n2843), .B(n4583), .Z(n3456) );
  HS65_LL_NOR2X2 U6137 ( .A(n4986), .B(n4583), .Z(n3552) );
  HS65_LL_NOR2X2 U6139 ( .A(n5320), .B(n4583), .Z(n4541) );
  HS65_LH_OAI22X1 U6140 ( .A(n4700), .B(n4583), .C(n3756), .D(n4701), .Z(n3595) );
  HS65_LL_OAI12X2 U6141 ( .A(n4583), .B(n4796), .C(n3518), .Z(n3520) );
  HS65_LL_OAI21X2 U6142 ( .A(n4583), .B(n4981), .C(n3718), .Z(n4494) );
  HS65_LL_NOR2X2 U6143 ( .A(n4700), .B(n4583), .Z(n3904) );
  HS65_LL_NOR2X2 U6145 ( .A(n4984), .B(n4583), .Z(n3840) );
  HS65_LH_NOR2X6 U6147 ( .A(n2854), .B(n4583), .Z(n3549) );
  HS65_LL_NAND2X7 U6150 ( .A(n3890), .B(n3889), .Z(n7867) );
  HS65_LH_OAI21X2 U6152 ( .A(n4293), .B(n4319), .C(n4292), .Z(n4294) );
  HS65_LL_AOI12X3 U6153 ( .A(n3803), .B(n3503), .C(n3502), .Z(n4319) );
  HS65_LH_OAI12X3 U6163 ( .A(n3802), .B(n3682), .C(n3684), .Z(n3502) );
  HS65_LL_OAI12X3 U6164 ( .A(n5209), .B(n3613), .C(n3615), .Z(n3803) );
  HS65_LL_NAND2X4 U6174 ( .A(n2881), .B(n6340), .Z(n6333) );
  HS65_LL_AOI12X2 U6179 ( .A(n4733), .B(n4732), .C(n4731), .Z(n4734) );
  HS65_LL_NOR3X2 U6190 ( .A(n4275), .B(n4274), .C(n4273), .Z(n4276) );
  HS65_LL_NAND2X2 U6196 ( .A(n5661), .B(n5660), .Z(n5662) );
  HS65_LH_NAND2X2 U6199 ( .A(n5618), .B(n5660), .Z(n4268) );
  HS65_LL_NOR3X1 U6202 ( .A(n4156), .B(n4153), .C(n4155), .Z(n4558) );
  HS65_LH_NOR2X2 U6203 ( .A(n5652), .B(n2893), .Z(n3823) );
  HS65_LL_NOR2X2 U6205 ( .A(n4465), .B(n4156), .Z(n3790) );
  HS65_LL_NOR2X2 U6208 ( .A(n4671), .B(n2893), .Z(n3955) );
  HS65_LL_IVX9 U6210 ( .A(n2893), .Z(n4544) );
  HS65_LL_OA12X9 U6213 ( .A(n5498), .B(n5497), .C(n5496), .Z(n5595) );
  HS65_LL_NOR2X2 U6215 ( .A(n8794), .B(n9049), .Z(\u_DataPath/cw_exmem_i [5])
         );
  HS65_LL_NAND2AX4 U6217 ( .A(n5640), .B(n5639), .Z(n5641) );
  HS65_LLS_XNOR2X3 U6219 ( .A(n2917), .B(n5637), .Z(n5638) );
  HS65_LL_NOR2X3 U6230 ( .A(n5397), .B(n4902), .Z(n3361) );
  HS65_LL_CNIVX3 U6234 ( .A(n5373), .Z(n3360) );
  HS65_LL_NAND2X4 U6235 ( .A(n5078), .B(n5077), .Z(n5079) );
  HS65_LH_IVX9 U6246 ( .A(\sub_x_53/A[17] ), .Z(n4984) );
  HS65_LH_NAND2X7 U6247 ( .A(n5667), .B(n4389), .Z(n4390) );
  HS65_LL_NAND3X3 U6249 ( .A(n3910), .B(n4022), .C(n3536), .Z(n4389) );
  HS65_LH_AOI12X3 U6257 ( .A(\sub_x_53/A[17] ), .B(n4588), .C(n3535), .Z(n3536) );
  HS65_LH_AOI12X3 U6262 ( .A(n4431), .B(n4349), .C(n4348), .Z(n4365) );
  HS65_LH_IVX9 U6265 ( .A(n9335), .Z(n9374) );
  HS65_LH_IVX9 U6266 ( .A(n9335), .Z(n9375) );
  HS65_LL_NOR2X2 U6269 ( .A(n4494), .B(n4500), .Z(n3905) );
  HS65_LH_AOI12X3 U6274 ( .A(n4516), .B(n4504), .C(n4503), .Z(n4510) );
  HS65_LL_NAND2X2 U6276 ( .A(\lte_x_59/B[18] ), .B(n4351), .Z(n3838) );
  HS65_LL_NOR2X2 U6277 ( .A(n4502), .B(n4501), .Z(n4503) );
  HS65_LH_NAND2X2 U6284 ( .A(n2858), .B(n4351), .Z(n4129) );
  HS65_LL_AOI211X1 U6285 ( .A(n2842), .B(n4351), .C(n4024), .D(n4023), .Z(
        n4579) );
  HS65_LH_NAND2X2 U6297 ( .A(\lte_x_59/B[9] ), .B(n4351), .Z(n4591) );
  HS65_LH_NAND2X2 U6298 ( .A(n2851), .B(n4351), .Z(n3543) );
  HS65_LH_NAND2X2 U6310 ( .A(\lte_x_59/B[16] ), .B(n4351), .Z(n3984) );
  HS65_LH_NAND2X2 U6311 ( .A(\lte_x_59/B[15] ), .B(n4351), .Z(n4059) );
  HS65_LL_NAND2X2 U6317 ( .A(\sub_x_53/A[25] ), .B(n4351), .Z(n3719) );
  HS65_LL_NAND2X4 U6332 ( .A(\lte_x_59/B[28] ), .B(n4351), .Z(n3759) );
  HS65_LH_OAI21X3 U6335 ( .A(n5394), .B(n5393), .C(n5392), .Z(n5414) );
  HS65_LL_NAND2X2 U6337 ( .A(n3327), .B(n9179), .Z(n3324) );
  HS65_LH_NAND2X2 U6338 ( .A(n3327), .B(n9343), .Z(n3157) );
  HS65_LL_NAND2X2 U6339 ( .A(n3327), .B(n9171), .Z(n3243) );
  HS65_LH_NAND2X2 U6347 ( .A(n3327), .B(n9342), .Z(n3148) );
  HS65_LH_NAND2X2 U6349 ( .A(n3327), .B(n9343), .Z(n3209) );
  HS65_LH_NAND2X2 U6355 ( .A(n3327), .B(n9342), .Z(n3172) );
  HS65_LH_NAND2X2 U6356 ( .A(n3327), .B(n9342), .Z(n3180) );
  HS65_LH_NAND2X2 U6360 ( .A(n3327), .B(n9185), .Z(n3263) );
  HS65_LH_NAND2X2 U6366 ( .A(n3327), .B(n9173), .Z(n3230) );
  HS65_LL_NAND2X2 U6367 ( .A(n3327), .B(n9175), .Z(n3328) );
  HS65_LH_NAND2X2 U6372 ( .A(n3327), .B(n9341), .Z(n3191) );
  HS65_LL_NAND2X4 U6392 ( .A(n3327), .B(n9033), .Z(n3314) );
  HS65_LL_NOR3X1 U6402 ( .A(n4471), .B(n4470), .C(n4469), .Z(n4472) );
  HS65_LL_OAI12X3 U6413 ( .A(n4468), .B(n5146), .C(n4467), .Z(n4469) );
  HS65_LH_AOI12X2 U6426 ( .A(n3474), .B(n4544), .C(n3868), .Z(n3869) );
  HS65_LL_NAND2AX4 U6435 ( .A(n5473), .B(n5472), .Z(n5481) );
  HS65_LL_NAND2X2 U6438 ( .A(n4805), .B(n4811), .Z(n5547) );
  HS65_LL_AOI12X2 U6447 ( .A(n5615), .B(n5248), .C(n5247), .Z(n5253) );
  HS65_LH_NOR2X2 U6450 ( .A(n4806), .B(n4506), .Z(n4505) );
  HS65_LH_NAND2X2 U6459 ( .A(n5448), .B(n4329), .Z(n4339) );
  HS65_LH_IVX2 U6460 ( .A(n4305), .Z(n4306) );
  HS65_LH_AOI12X6 U6474 ( .A(n4303), .B(n4305), .C(n4231), .Z(n4235) );
  HS65_LL_OAI12X2 U6480 ( .A(n4331), .B(n4328), .C(n5448), .Z(n5452) );
  HS65_LL_OAI12X2 U6490 ( .A(n4331), .B(n4328), .C(n5448), .Z(n4305) );
  HS65_LL_NAND2X4 U6493 ( .A(n9369), .B(n9042), .Z(n8294) );
  HS65_LL_IVX4 U6496 ( .A(\u_DataPath/dataOut_exe_i [29]), .Z(n4213) );
  HS65_LL_NAND2X2 U6501 ( .A(n9366), .B(n9079), .Z(n8312) );
  HS65_LL_NAND2X2 U6504 ( .A(n9368), .B(n9006), .Z(n8432) );
  HS65_LL_NAND2X4 U6507 ( .A(n9368), .B(n9101), .Z(n8398) );
  HS65_LL_NAND2X4 U6519 ( .A(n9366), .B(n9043), .Z(n7836) );
  HS65_LL_NAND2X4 U6530 ( .A(n9365), .B(n9044), .Z(n8290) );
  HS65_LL_NAND2X4 U6531 ( .A(n9366), .B(n9015), .Z(n8340) );
  HS65_LL_NAND2X4 U6532 ( .A(n8166), .B(n6138), .Z(n6149) );
  HS65_LL_AOI22X3 U6538 ( .A(n8868), .B(n9034), .C(n9368), .D(n8946), .Z(n7851) );
  HS65_LL_NAND2X2 U6539 ( .A(n9369), .B(n9014), .Z(n8307) );
  HS65_LL_NAND2X2 U6547 ( .A(n9365), .B(n9249), .Z(n8436) );
  HS65_LL_NAND2X2 U6551 ( .A(n9369), .B(n9045), .Z(n8333) );
  HS65_LL_NAND2X4 U6554 ( .A(n4322), .B(n5210), .Z(n4324) );
  HS65_LL_AOI21X2 U6556 ( .A(n4322), .B(n5211), .C(n4321), .Z(n4323) );
  HS65_LL_NOR2X6 U6557 ( .A(n3682), .B(n3800), .Z(n3503) );
  HS65_LL_NOR2X5 U6558 ( .A(n2853), .B(n5567), .Z(n3800) );
  HS65_LL_NAND2X11 U6560 ( .A(n3157), .B(n3156), .Z(n5567) );
  HS65_LL_NOR3X4 U6565 ( .A(n5486), .B(n5485), .C(n5484), .Z(n5487) );
  HS65_LL_CBI4I1X3 U6567 ( .A(n5508), .B(n5367), .C(n5366), .D(n5365), .Z(
        n5484) );
  HS65_LL_AOI12X2 U6568 ( .A(n5643), .B(n5155), .C(n5154), .Z(n5156) );
  HS65_LL_OAI12X2 U6572 ( .A(n5153), .B(n5152), .C(n5151), .Z(n5154) );
  HS65_LL_IVX7 U6585 ( .A(n5646), .Z(n5229) );
  HS65_LL_NOR2X2 U6591 ( .A(\lte_x_59/B[3] ), .B(n5089), .Z(n4570) );
  HS65_LL_AOI12X2 U6594 ( .A(n4638), .B(n4645), .C(n4640), .Z(n4145) );
  HS65_LL_CNIVX3 U6595 ( .A(n9376), .Z(n3327) );
  HS65_LL_CNIVX3 U6598 ( .A(n3593), .Z(n5425) );
  HS65_LL_AND2X4 U6603 ( .A(n3132), .B(n7802), .Z(n3133) );
  HS65_LL_AOI21X2 U6605 ( .A(n5229), .B(n3723), .C(n3722), .Z(n3724) );
  HS65_LL_AOI12X2 U6618 ( .A(n3727), .B(n5624), .C(n3726), .Z(n3728) );
  HS65_LH_OAI21X2 U6619 ( .A(n3725), .B(n5656), .C(n3724), .Z(n3726) );
  HS65_LL_MUXI21X5 U6620 ( .D0(n2972), .D1(n2971), .S0(
        \u_DataPath/cw_towb_i [0]), .Z(n8393) );
  HS65_LL_CNIVX3 U6623 ( .A(\u_DataPath/from_mem_data_out_i [4]), .Z(n2971) );
  HS65_LL_NAND3X2 U6624 ( .A(n4163), .B(n4162), .C(n4161), .Z(n5671) );
  HS65_LL_NAND2X5 U6625 ( .A(n8177), .B(n7802), .Z(n8486) );
  HS65_LL_IVX7 U6626 ( .A(n4953), .Z(n4148) );
  HS65_LH_AOI12X2 U6628 ( .A(n5144), .B(n4875), .C(n4118), .Z(n4125) );
  HS65_LL_IVX4 U6632 ( .A(n4113), .Z(n4875) );
  HS65_LH_OAI21X2 U6636 ( .A(n5173), .B(n4117), .C(n4116), .Z(n4118) );
  HS65_LL_AOI21X2 U6637 ( .A(n3529), .B(n4114), .C(n5041), .Z(n4115) );
  HS65_LL_NAND2X2 U6638 ( .A(n5648), .B(n5040), .Z(n4114) );
  HS65_LL_OAI21X3 U6652 ( .A(n4821), .B(n4817), .C(n4819), .Z(n4538) );
  HS65_LL_NAND2X4 U6654 ( .A(\lte_x_59/B[1] ), .B(n3294), .Z(n4819) );
  HS65_LL_NOR2X5 U6657 ( .A(\lte_x_59/B[1] ), .B(n3294), .Z(n4817) );
  HS65_LH_IVX2 U6658 ( .A(n4805), .Z(n3294) );
  HS65_LL_AOI21X4 U6659 ( .A(n5624), .B(n4446), .C(n4445), .Z(n4447) );
  HS65_LL_NAND3X5 U6661 ( .A(n4444), .B(n4443), .C(n4442), .Z(n4445) );
  HS65_LH_NOR2X2 U6662 ( .A(n4855), .B(n4435), .Z(n4436) );
  HS65_LL_AND2ABX9 U6663 ( .A(n4458), .B(n4842), .Z(n5618) );
  HS65_LL_NOR3X7 U6664 ( .A(n4782), .B(n4783), .C(n4784), .Z(n4785) );
  HS65_LL_NAND3X3 U6666 ( .A(n5516), .B(n5517), .C(n5408), .Z(n4684) );
  HS65_LL_NOR2X5 U6667 ( .A(n5406), .B(n5294), .Z(n5408) );
  HS65_LL_OAI112X1 U6670 ( .A(n9129), .B(n8880), .C(n8308), .D(n9086), .Z(
        \u_DataPath/from_mem_data_out_i [15]) );
  HS65_LLS_XOR2X3 U6671 ( .A(n4635), .B(n4634), .Z(n4636) );
  HS65_LL_AOI12X2 U6675 ( .A(n4633), .B(n4632), .C(n4631), .Z(n4634) );
  HS65_LL_AOI12X12 U6687 ( .A(n5906), .B(n5908), .C(n5740), .Z(n5746) );
  HS65_LL_OAI12X2 U6701 ( .A(n5855), .B(n5854), .C(n5853), .Z(n5856) );
  HS65_LH_OAI21X3 U6704 ( .A(n5867), .B(n5817), .C(n5819), .Z(n5813) );
  HS65_LL_NOR2X3 U6705 ( .A(n3629), .B(n3747), .Z(n5446) );
  HS65_LL_NOR2AX3 U6706 ( .A(n4233), .B(n4332), .Z(n4234) );
  HS65_LH_OAI21X2 U6707 ( .A(n3747), .B(n3632), .C(n3749), .Z(n3633) );
  HS65_LH_OAI12X2 U6708 ( .A(n4333), .B(n4332), .C(n4331), .Z(n4334) );
  HS65_LL_NOR2X6 U6710 ( .A(n2853), .B(n3384), .Z(n3747) );
  HS65_LL_NAND2AX7 U6714 ( .A(n7634), .B(n7622), .Z(n4227) );
  HS65_LL_NAND2AX4 U6718 ( .A(n7634), .B(n4380), .Z(n4416) );
  HS65_LL_AND2X4 U6719 ( .A(n5217), .B(n4301), .Z(n5708) );
  HS65_LL_NAND2X2 U6721 ( .A(n5217), .B(n3510), .Z(n3511) );
  HS65_LL_AND2X4 U6734 ( .A(n5217), .B(n3849), .Z(n3850) );
  HS65_LL_NAND2X2 U6741 ( .A(n5217), .B(n3944), .Z(n3945) );
  HS65_LL_NAND2X4 U6745 ( .A(n5217), .B(n3995), .Z(n3996) );
  HS65_LH_NAND2X2 U6753 ( .A(n5217), .B(n4479), .Z(n4485) );
  HS65_LL_IVX9 U6768 ( .A(n7634), .Z(n5643) );
  HS65_LL_CNIVX3 U6778 ( .A(n5217), .Z(n7634) );
  HS65_LH_NAND2X2 U6796 ( .A(\u_DataPath/cw_to_ex_i [3]), .B(n5492), .Z(n3450)
         );
  HS65_LL_NOR2X2 U6797 ( .A(\u_DataPath/cw_to_ex_i [3]), .B(
        \u_DataPath/cw_to_ex_i [4]), .Z(n3470) );
  HS65_LL_NAND2X5 U6799 ( .A(n7631), .B(n5280), .Z(n5281) );
  HS65_LLS_XNOR2X6 U6800 ( .A(n5279), .B(n5278), .Z(n5280) );
  HS65_LL_MX41X4 U6801 ( .D0(n8440), .S0(n9289), .D1(n8441), .S1(n9274), .D2(
        n8439), .S2(n9296), .D3(n8438), .S3(n9281), .Z(
        \u_DataPath/from_mem_data_out_i [0]) );
  HS65_LL_OAI21X2 U6804 ( .A(n4534), .B(n4533), .C(n2928), .Z(n5705) );
  HS65_LL_NOR3X4 U6812 ( .A(n4532), .B(n4531), .C(n4530), .Z(n2928) );
  HS65_LH_IVX9 U6813 ( .A(\u_DataPath/from_mem_data_out_i [0]), .Z(n3015) );
  HS65_LL_NOR2X2 U6819 ( .A(n4700), .B(n5129), .Z(n3779) );
  HS65_LL_NAND2X7 U6840 ( .A(\lte_x_59/B[15] ), .B(n4677), .Z(n3893) );
  HS65_LH_CNIVX7 U6850 ( .A(n5062), .Z(n4677) );
  HS65_LL_NAND3X2 U6851 ( .A(n8775), .B(n9169), .C(n8078), .Z(n8079) );
  HS65_LL_NOR2X9 U6867 ( .A(\u_DataPath/cw_to_ex_i [4]), .B(n5120), .Z(n3422)
         );
  HS65_LH_IVX9 U6868 ( .A(n3422), .Z(n3423) );
  HS65_LL_NAND2X4 U6870 ( .A(n5491), .B(n3422), .Z(n3442) );
  HS65_LL_NAND3X2 U6916 ( .A(n5090), .B(n5474), .C(n5319), .Z(n4662) );
  HS65_LL_NOR2X3 U6923 ( .A(n4661), .B(n5548), .Z(n5319) );
  HS65_LL_NAND2X5 U6927 ( .A(\sub_x_53/A[2] ), .B(n3415), .Z(n4573) );
  HS65_LL_OAI12X2 U6928 ( .A(n5546), .B(n5318), .C(n4662), .Z(n4669) );
  HS65_LL_NAND2X2 U6931 ( .A(n5090), .B(n4573), .Z(n5546) );
  HS65_LL_IVX7 U6943 ( .A(\u_DataPath/from_mem_data_out_i [2]), .Z(n2933) );
  HS65_LL_NAND2X7 U6957 ( .A(n3512), .B(n3511), .Z(n3513) );
  HS65_LLS_XNOR2X6 U6963 ( .A(n3509), .B(n3508), .Z(n3510) );
  HS65_LL_IVX7 U6964 ( .A(\u_DataPath/from_mem_data_out_i [3]), .Z(n2969) );
  HS65_LL_OAI22X1 U6971 ( .A(n3333), .B(\u_DataPath/dataOut_exe_i [5]), .C(
        n8391), .D(n3340), .Z(n3334) );
  HS65_LH_NOR2X5 U6975 ( .A(n8391), .B(n9401), .Z(n4654) );
  HS65_LLS_XNOR2X3 U6984 ( .A(n4884), .B(n4883), .Z(n4885) );
  HS65_LL_NOR3X4 U6988 ( .A(n3465), .B(n3464), .C(n3463), .Z(n3466) );
  HS65_LL_NAND2AX4 U7002 ( .A(n3438), .B(n3437), .Z(n3465) );
  HS65_LL_OAI31X2 U7006 ( .A(n5177), .B(n4581), .C(n3713), .D(n3454), .Z(n3464) );
  HS65_LH_NAND2X5 U7010 ( .A(n5170), .B(n5667), .Z(n3437) );
  HS65_LL_NOR3X4 U7012 ( .A(\u_DataPath/u_idexreg/N15 ), .B(n8103), .C(
        \u_DataPath/u_idexreg/N10 ), .Z(n8126) );
  HS65_LH_NAND2X7 U7014 ( .A(n7631), .B(n4414), .Z(n4415) );
  HS65_LL_NOR2X3 U7015 ( .A(\lte_x_59/B[6] ), .B(n2865), .Z(n4643) );
  HS65_LL_NAND2X4 U7037 ( .A(n3323), .B(n3322), .Z(n3325) );
  HS65_LL_NAND3X5 U7045 ( .A(n5220), .B(n5219), .C(n5218), .Z(n5221) );
  HS65_LL_NAND2X4 U7048 ( .A(n5217), .B(n5216), .Z(n5218) );
  HS65_LL_NOR2X5 U7049 ( .A(\lte_x_59/B[16] ), .B(n5021), .Z(n3560) );
  HS65_LL_NAND2X5 U7051 ( .A(n3207), .B(n8526), .Z(n3208) );
  HS65_LLS_XNOR2X3 U7063 ( .A(n5215), .B(n5214), .Z(n5216) );
  HS65_LL_NAND2X4 U7069 ( .A(n5672), .B(n6122), .Z(n4277) );
  HS65_LL_NAND3X5 U7082 ( .A(n4266), .B(n4265), .C(n4264), .Z(n6122) );
  HS65_LL_AND2X4 U7085 ( .A(n9211), .B(n9366), .Z(n8424) );
  HS65_LL_CNIVX7 U7097 ( .A(\u_DataPath/dataOut_exe_i [1]), .Z(n8177) );
  HS65_LL_NOR2X3 U7098 ( .A(n4701), .B(n4582), .Z(n3953) );
  HS65_LL_NAND2X7 U7100 ( .A(n8166), .B(n6145), .Z(n6152) );
  HS65_LH_IVX2 U7104 ( .A(\u_DataPath/jaddr_i [25]), .Z(n8166) );
  HS65_LL_AND2ABX18 U7109 ( .A(n3425), .B(n5088), .Z(n4836) );
  HS65_LL_AOI21X2 U7114 ( .A(n5661), .B(n5239), .C(n5238), .Z(n5245) );
  HS65_LL_IVX7 U7121 ( .A(n4609), .Z(n5239) );
  HS65_LL_AOI21X2 U7154 ( .A(n5229), .B(n5228), .C(n5227), .Z(n5246) );
  HS65_LL_NAND3AX6 U7160 ( .A(n3829), .B(n3828), .C(n3827), .Z(n3844) );
  HS65_LL_CNIVX3 U7161 ( .A(n4840), .Z(n3858) );
  HS65_LL_NOR2AX3 U7172 ( .A(n3789), .B(n2860), .Z(n3820) );
  HS65_LLS_XNOR2X3 U7173 ( .A(n4482), .B(n4645), .Z(n4483) );
  HS65_LL_AOI21X2 U7180 ( .A(n4646), .B(n4645), .C(n4644), .Z(n4647) );
  HS65_LL_OAI21X2 U7183 ( .A(n3394), .B(n8485), .C(n3395), .Z(n3293) );
  HS65_LL_MX41X4 U7194 ( .D0(n8441), .S0(n9275), .D1(n8440), .S1(n9290), .D2(
        n9297), .S2(n8439), .D3(n8438), .S3(n9282), .Z(
        \u_DataPath/from_mem_data_out_i [1]) );
  HS65_LL_NAND4ABX3 U7197 ( .A(n8106), .B(n8105), .C(n8104), .D(n8126), .Z(
        \u_DataPath/cw_to_ex_i [2]) );
  HS65_LL_NAND2X2 U7208 ( .A(n5667), .B(n3522), .Z(n3523) );
  HS65_LL_NOR2X2 U7210 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5079), .Z(n5117)
         );
  HS65_LH_OAI21X2 U7217 ( .A(n5173), .B(n5204), .C(n3880), .Z(n3881) );
  HS65_LH_AOI22X1 U7218 ( .A(n4951), .B(n4615), .C(n5667), .D(n4614), .Z(n4619) );
  HS65_LH_NAND2X2 U7223 ( .A(n5667), .B(n5228), .Z(n3714) );
  HS65_LL_NOR2X2 U7224 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5119), .Z(n4782)
         );
  HS65_LL_NAND2X2 U7225 ( .A(n5667), .B(n5174), .Z(n4848) );
  HS65_LH_NOR2X2 U7233 ( .A(n5173), .B(n4357), .Z(n4358) );
  HS65_LL_OAI21X2 U7245 ( .A(n5173), .B(n4526), .C(n4525), .Z(n4531) );
  HS65_LL_NAND2X2 U7255 ( .A(n5667), .B(n5617), .Z(n4267) );
  HS65_LH_OAI22X1 U7275 ( .A(n4435), .B(n5173), .C(n4954), .D(n3858), .Z(n3829) );
  HS65_LL_NOR2X2 U7285 ( .A(n5173), .B(n4355), .Z(n3597) );
  HS65_LL_AOI12X2 U7306 ( .A(n5667), .B(n5243), .C(n5242), .Z(n5244) );
  HS65_LL_NAND2X2 U7308 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(
        \u_DataPath/cw_to_ex_i [2]), .Z(n4965) );
  HS65_LL_NOR2X2 U7314 ( .A(\u_DataPath/u_idexreg/N3 ), .B(n5463), .Z(n5469)
         );
  HS65_LL_NOR2X2 U7333 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n7617), .Z(n5217)
         );
  HS65_LL_NAND2X4 U7356 ( .A(n5463), .B(n5492), .Z(n5120) );
  HS65_LL_NAND2X4 U7376 ( .A(\u_DataPath/cw_to_ex_i [1]), .B(n5492), .Z(n3417)
         );
  HS65_LL_IVX2 U7379 ( .A(\u_DataPath/cw_to_ex_i [1]), .Z(n5463) );
  HS65_LH_IVX2 U7381 ( .A(n8704), .Z(n3122) );
  HS65_LL_AND3X18 U7386 ( .A(n8101), .B(n8072), .C(n8071), .Z(n9376) );
  HS65_LL_OA12X4 U7387 ( .A(n9242), .B(n8453), .C(n7913), .Z(n9377) );
  HS65_LH_OA222X4 U7393 ( .A(n9166), .B(n8898), .C(n9051), .D(n9127), .E(n8880), .F(n9268), .Z(n9378) );
  HS65_LL_OA12X4 U7394 ( .A(n9268), .B(n8453), .C(n7913), .Z(n9379) );
  HS65_LL_OA12X4 U7395 ( .A(n9123), .B(n8453), .C(n7913), .Z(n9380) );
  HS65_LH_IVX2 U7396 ( .A(n8267), .Z(\u_DataPath/dataOut_exe_i [8]) );
  HS65_LL_OA112X4 U7397 ( .A(n9246), .B(n8880), .C(n8291), .D(n9086), .Z(n9381) );
  HS65_LL_OA12X4 U7399 ( .A(n9120), .B(n8453), .C(n9086), .Z(n9383) );
  HS65_LL_OA12X4 U7401 ( .A(n9247), .B(n8453), .C(n9086), .Z(n9384) );
  HS65_LL_OA12X4 U7404 ( .A(n9121), .B(n8453), .C(n7913), .Z(n9385) );
  HS65_LL_OA112X4 U7405 ( .A(n9244), .B(n8880), .C(n8346), .D(n9086), .Z(n9386) );
  HS65_LL_OA12X4 U7408 ( .A(n9124), .B(n8453), .C(n7913), .Z(n9387) );
  HS65_LL_OA12X4 U7409 ( .A(n9243), .B(n8453), .C(n9086), .Z(n9388) );
  HS65_LH_OA12X9 U7411 ( .A(n9245), .B(n8453), .C(n7913), .Z(n9389) );
  HS65_LL_OA12X4 U7413 ( .A(n9125), .B(n8453), .C(n7913), .Z(n9391) );
  HS65_LL_OA12X4 U7414 ( .A(n9248), .B(n8453), .C(n7913), .Z(n9392) );
  HS65_LL_OA12X4 U7415 ( .A(n9244), .B(n8453), .C(n7913), .Z(n9393) );
  HS65_LL_OA12X4 U7450 ( .A(n9126), .B(n8453), .C(n7913), .Z(n9394) );
  HS65_LL_OA12X4 U7454 ( .A(n9129), .B(n8453), .C(n9086), .Z(n9395) );
  HS65_LL_OA112X4 U7456 ( .A(n8880), .B(n9245), .C(n8273), .D(n9086), .Z(n9396) );
  HS65_LH_IVX2 U7461 ( .A(n8297), .Z(\u_DataPath/dataOut_exe_i [7]) );
  HS65_LL_OA112X4 U7466 ( .A(n9247), .B(n8880), .C(n8341), .D(n9086), .Z(n9397) );
  HS65_LL_OA112X4 U7473 ( .A(n9242), .B(n8880), .C(n8334), .D(n9086), .Z(n9398) );
  HS65_LH_OA22X4 U7480 ( .A(n8906), .B(n9269), .C(n9140), .D(n8758), .Z(n9399)
         );
  HS65_LH_OA22X4 U7494 ( .A(n8906), .B(n9270), .C(n9140), .D(n8760), .Z(n9400)
         );
  HS65_LL_OR3ABCX35 U7500 ( .A(n3217), .B(n2966), .C(n3216), .Z(n9401) );
  HS65_LH_IVX18 U7524 ( .A(n2846), .Z(n2847) );
  HS65_LLS_XNOR2X3 U7531 ( .A(n4821), .B(n4820), .Z(n9402) );
  HS65_LH_AO22X4 U7551 ( .A(n9261), .B(n9136), .C(n9134), .D(n8936), .Z(n9403)
         );
  HS65_LH_AO22X4 U7555 ( .A(n9056), .B(n9136), .C(n9134), .D(n8956), .Z(n9404)
         );
  HS65_LH_AO22X4 U7575 ( .A(n9089), .B(n9136), .C(n9134), .D(n8953), .Z(n9405)
         );
  HS65_LH_AO22X4 U7577 ( .A(n9094), .B(n9136), .C(n9134), .D(n8957), .Z(n9406)
         );
  HS65_LH_AO22X4 U7583 ( .A(n9259), .B(n9136), .C(n9134), .D(n8950), .Z(n9407)
         );
  HS65_LH_AO22X4 U7584 ( .A(n9091), .B(n9136), .C(n9134), .D(n8955), .Z(n9408)
         );
  HS65_LH_AO22X4 U7591 ( .A(n8881), .B(n9136), .C(n9134), .D(n8954), .Z(n9409)
         );
  HS65_LH_AO22X4 U7598 ( .A(n9095), .B(n9136), .C(n9134), .D(n8959), .Z(n9410)
         );
  HS65_LH_AO22X4 U7599 ( .A(n9106), .B(n9136), .C(n9134), .D(n8958), .Z(n9411)
         );
  HS65_LH_AO22X4 U7604 ( .A(n9088), .B(n9136), .C(n9134), .D(n9064), .Z(n9412)
         );
  HS65_LH_AO22X4 U7605 ( .A(n9096), .B(n9136), .C(n9134), .D(n8952), .Z(n9413)
         );
  HS65_LH_AO22X4 U7606 ( .A(n9071), .B(n9136), .C(n9133), .D(n8977), .Z(n9414)
         );
  HS65_LH_AO22X4 U7660 ( .A(n9271), .B(n9188), .C(n9133), .D(n8990), .Z(n9415)
         );
  HS65_LH_AO22X4 U7676 ( .A(n9257), .B(n9188), .C(n9133), .D(n9023), .Z(n9416)
         );
  HS65_LH_AO22X4 U7677 ( .A(n9107), .B(n9188), .C(n9133), .D(n9024), .Z(n9417)
         );
  HS65_LH_AO22X4 U7686 ( .A(n9136), .B(n9200), .C(n9134), .D(n8949), .Z(n9418)
         );
  HS65_LH_IVX7 U7710 ( .A(n8704), .Z(n2784) );
  HS65_LH_AO22X4 U7727 ( .A(n9192), .B(n9265), .C(n9132), .D(n9067), .Z(n9419)
         );
  HS65_LH_AO22X4 U7734 ( .A(n9192), .B(n9161), .C(n9132), .D(n8989), .Z(n9420)
         );
  HS65_LH_AO22X4 U7743 ( .A(n9192), .B(n9143), .C(n9132), .D(n8995), .Z(n9421)
         );
  HS65_LH_AO22X4 U7746 ( .A(n9192), .B(n9158), .C(n9132), .D(n8978), .Z(n9422)
         );
  HS65_LH_AO22X4 U7749 ( .A(n9192), .B(n9157), .C(n9132), .D(n8973), .Z(n9423)
         );
  HS65_LH_AO22X4 U7751 ( .A(n9192), .B(n9162), .C(n9132), .D(n8986), .Z(n9424)
         );
  HS65_LH_AO22X4 U7763 ( .A(n9192), .B(n9160), .C(n9132), .D(n9087), .Z(n9425)
         );
  HS65_LH_AO22X4 U7764 ( .A(n9192), .B(n9156), .C(n9132), .D(n8962), .Z(n9426)
         );
  HS65_LH_AO22X4 U7771 ( .A(n9192), .B(n9155), .C(n9132), .D(n8976), .Z(n9427)
         );
  HS65_LH_AO22X4 U7776 ( .A(n9191), .B(n9163), .C(n9131), .D(n8991), .Z(n9428)
         );
  HS65_LH_AO22X4 U7779 ( .A(n9191), .B(n9159), .C(n9131), .D(n8988), .Z(n9429)
         );
  HS65_LH_NOR2X2 U7780 ( .A(n9233), .B(n7117), .Z(n2877) );
  HS65_LH_NAND4ABX3 U7809 ( .A(n9347), .B(n8755), .C(n9016), .D(n8071), .Z(
        \u_DataPath/cw_exmem_i [10]) );
  HS65_LL_DFPQX9 clk_r_REG490_S3 ( .D(n8635), .CP(clk), .Q(n9066) );
  HS65_LL_OAI211X5 U3847 ( .A(n9149), .B(n9012), .C(n8877), .D(n8093), .Z(
        \u_DataPath/cw_to_ex_i [3]) );
  HS65_LL_NAND2AX7 U6275 ( .A(n4867), .B(n4866), .Z(n5686) );
  HS65_LH_DFPQX4 clk_r_REG48_S1 ( .D(n8580), .CP(clk), .Q(n3023) );
  HS65_LH_DFPQX4 clk_r_REG435_S3 ( .D(n8270), .CP(clk), .Q(n9081) );
  HS65_LL_DFPQX4 clk_r_REG387_S2 ( .D(\u_DataPath/data_read_ex_2_i [0]), .CP(
        clk), .Q(n9431) );
  HS65_LH_DFPQX4 clk_r_REG431_S2 ( .D(n9115), .CP(clk), .Q(n9114) );
  HS65_LL_DFPQNX9 clk_r_REG450_S1 ( .D(n8137), .CP(clk), .QN(
        \u_DataPath/cw_towb_i [0]) );
  HS65_LH_DFPQX9 clk_r_REG76_S2 ( .D(n8473), .CP(clk), .Q(n9027) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[31][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N92 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[18][24]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N137 ), .D(n7984), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][24] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[26][27]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N129 ), .D(n7926), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7986), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][9]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n8013), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][9] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[30][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N125 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[30][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][0]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7998), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][0] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[29][17]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N126 ), .D(n7987), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[29][17] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][22]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7977), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][22] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][21]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7965), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][21] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][23]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7995), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][23] ) );
  HS65_LH_LDHQX4 \u_DataPath/u_decode_unit/reg_file0/bank_register_reg[28][11]  ( 
        .G(\u_DataPath/u_decode_unit/reg_file0/N127 ), .D(n7941), .Q(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[28][11] ) );
  HS65_LH_DFPQX4 clk_r_REG660_S1 ( .D(Data_out_fromRAM[24]), .CP(clk), .Q(
        n9296) );
  HS65_LH_DFPQX4 clk_r_REG686_S1 ( .D(Data_out_fromRAM[6]), .CP(clk), .Q(n9280) );
  HS65_LH_DFPQX4 clk_r_REG395_S2 ( .D(n2851), .CP(clk), .Q(n9261) );
  HS65_LH_DFPQX9 clk_r_REG657_S1 ( .D(n8319), .CP(clk), .Q(n9243) );
  HS65_LH_DFPQX4 clk_r_REG368_S2 ( .D(n9212), .CP(clk), .Q(n9211) );
  HS65_LH_DFPQX4 clk_r_REG270_S1 ( .D(\u_DataPath/branch_target_i [9]), .CP(
        clk), .Q(n9195) );
  HS65_LH_DFPQX4 clk_r_REG589_S2 ( .D(n9179), .CP(clk), .Q(n9178) );
  HS65_LH_DFPRQX4 clk_r_REG512_S1 ( .D(n7897), .CP(clk), .RN(n7879), .Q(n9132)
         );
  HS65_LH_DFPQX4 clk_r_REG451_S1 ( .D(\u_DataPath/cw_tomem_i [4]), .CP(clk), 
        .Q(n9112) );
  HS65_LH_DFPQX4 clk_r_REG60_S5 ( .D(\lte_x_59/B[6] ), .CP(clk), .Q(n9095) );
  HS65_LH_DFPQX4 clk_r_REG149_S2 ( .D(\u_DataPath/u_execute/link_value_i [28]), 
        .CP(clk), .Q(n9057) );
  HS65_LH_DFPQX4 clk_r_REG121_S2 ( .D(\u_DataPath/u_execute/link_value_i [10]), 
        .CP(clk), .Q(n9042) );
  HS65_LH_DFPQX4 clk_r_REG573_S3 ( .D(n8086), .CP(clk), .Q(n9007) );
  HS65_LH_DFPRQX4 clk_r_REG154_S4 ( .D(\u_DataPath/pc_4_i [22]), .CP(clk), 
        .RN(n9354), .Q(n8988) );
  HS65_LH_DFPQX4 clk_r_REG268_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [11]), 
        .CP(clk), .Q(n8950) );
  HS65_LH_DFPQX4 clk_r_REG378_S2 ( .D(\u_DataPath/u_execute/resAdd1_i [1]), 
        .CP(clk), .Q(n8935) );
  HS65_LH_DFPQX4 clk_r_REG122_S1 ( .D(\u_DataPath/branch_target_i [13]), .CP(
        clk), .Q(n8919) );
  HS65_LH_DFPQX4 clk_r_REG61_S5 ( .D(n8479), .CP(clk), .Q(n8901) );
  HS65_LH_DFPQX4 clk_r_REG146_S2 ( .D(\u_DataPath/u_execute/link_value_i [29]), 
        .CP(clk), .Q(n8870) );
  HS65_LH_DFPRQX4 clk_r_REG604_S3 ( .D(\u_DataPath/immediate_ext_dec_i [13]), 
        .CP(clk), .RN(n9354), .Q(n8790) );
  HS65_LH_DFPRQX4 clk_r_REG559_S3 ( .D(\u_DataPath/jaddr_i [22]), .CP(clk), 
        .RN(n9354), .Q(n8765) );
  HS65_LH_DFPQX4 clk_r_REG29_S2 ( .D(\u_DataPath/mem_writedata_out_i [27]), 
        .CP(clk), .Q(n8748) );
  HS65_LH_DFPQX4 clk_r_REG81_S1 ( .D(\u_DataPath/mem_writedata_out_i [24]), 
        .CP(clk), .Q(n8732) );
  HS65_LL_IVX9 U3856 ( .A(n8898), .Z(n8399) );
  HS65_LL_NAND2X7 U7793 ( .A(n9102), .B(n9066), .Z(n8114) );
  HS65_LH_OAI12X3 U6125 ( .A(n9190), .B(n9027), .C(n8307), .Z(
        \u_DataPath/dataOut_exe_i [15]) );
  HS65_LL_BFX18 U4321 ( .A(n9401), .Z(n7868) );
  HS65_LL_NOR2X6 U3948 ( .A(n3214), .B(n3213), .Z(\lte_x_59/B[8] ) );
  HS65_LL_OAI12X3 U3808 ( .A(n3349), .B(n4712), .C(n3348), .Z(n3419) );
  HS65_LH_IVX9 U6106 ( .A(n5053), .Z(n2871) );
  HS65_LL_OAI12X6 U6982 ( .A(n4654), .B(n3339), .C(n4655), .Z(n5040) );
  HS65_LL_AOI21X2 U6075 ( .A(n9376), .B(n7846), .C(n3419), .Z(n3430) );
  HS65_LL_NOR3AX9 U3639 ( .A(n4971), .B(n4973), .C(n3059), .Z(\lte_x_59/B[28] ) );
  HS65_LL_NOR2X6 U5623 ( .A(n3086), .B(n3085), .Z(\lte_x_59/B[18] ) );
  HS65_LL_AND2ABX18 U3927 ( .A(n3096), .B(n3095), .Z(\lte_x_59/B[16] ) );
  HS65_LL_NAND2X7 U5585 ( .A(n3421), .B(n3422), .Z(n5179) );
  HS65_LL_IVX9 U3750 ( .A(n3443), .Z(n3529) );
  HS65_LL_IVX27 U3472 ( .A(n4795), .Z(n2864) );
  HS65_LH_IVX9 U6673 ( .A(n5180), .Z(n3382) );
  HS65_LH_NOR2AX6 U3718 ( .A(n3967), .B(n2872), .Z(n4550) );
  HS65_LL_NOR2AX6 U3894 ( .A(n3210), .B(n4420), .Z(n5194) );
  HS65_LH_NOR2AX3 U3700 ( .A(n9019), .B(n2994), .Z(n3014) );
  HS65_LL_IVX18 U3452 ( .A(n2774), .Z(Data_in[23]) );
  HS65_LL_IVX18 U3453 ( .A(n2776), .Z(Data_in[9]) );
  HS65_LL_IVX18 U3454 ( .A(n2778), .Z(Data_in[18]) );
  HS65_LL_IVX18 U3459 ( .A(n2819), .Z(Data_in[22]) );
  HS65_LL_IVX18 U3460 ( .A(n2821), .Z(Data_in[13]) );
  HS65_LL_IVX18 U3461 ( .A(n2838), .Z(Data_in[19]) );
  HS65_LL_CNBFX14 U3699 ( .A(n3014), .Z(Data_in[8]) );
  HS65_LL_IVX18 U3439 ( .A(n2787), .Z(Address_toRAM[21]) );
  HS65_LL_IVX18 U3440 ( .A(n2789), .Z(Address_toRAM[20]) );
  HS65_LL_IVX18 U3441 ( .A(n2791), .Z(Address_toRAM[23]) );
  HS65_LL_IVX18 U3442 ( .A(n2793), .Z(Address_toRAM[22]) );
  HS65_LL_IVX18 U3443 ( .A(n2795), .Z(Address_toRAM[19]) );
  HS65_LL_IVX18 U3444 ( .A(n2797), .Z(Address_toRAM[18]) );
  HS65_LL_IVX18 U3445 ( .A(n2799), .Z(Address_toRAM[28]) );
  HS65_LL_IVX18 U3450 ( .A(n2801), .Z(Address_toRAM[27]) );
  HS65_LL_IVX18 U3456 ( .A(n2805), .Z(Address_toRAM[6]) );
  HS65_LL_IVX18 U3458 ( .A(n2809), .Z(Address_toRAM[9]) );
  HS65_LL_IVX18 U3451 ( .A(n2811), .Z(Data_in[27]) );
  HS65_LL_IVX18 U3524 ( .A(n2815), .Z(Data_in[29]) );
  HS65_LL_IVX18 U3525 ( .A(n2813), .Z(Data_in[28]) );
  HS65_LL_IVX18 U3527 ( .A(n2817), .Z(Data_in[30]) );
  HS65_LL_IVX18 U3455 ( .A(n2803), .Z(Address_toRAM[10]) );
  HS65_LL_IVX18 U3457 ( .A(n2807), .Z(Address_toRAM[8]) );
  HS65_LL_IVX18 U3449 ( .A(n2784), .Z(addr_to_iram[14]) );
  HS65_LL_NAND2X7 U6252 ( .A(n3395), .B(n3394), .Z(n3396) );
  HS65_LH_BFX35 U3435 ( .A(n2986), .Z(n3116) );
  HS65_LL_IVX18 U3436 ( .A(n3120), .Z(addr_to_iram[23]) );
  HS65_LL_IVX18 U3510 ( .A(n7785), .Z(addr_to_iram[28]) );
  HS65_LL_IVX18 U3513 ( .A(n3121), .Z(addr_to_iram[22]) );
  HS65_LH_BFX9 U3514 ( .A(n2994), .Z(n3115) );
  HS65_LL_NAND2X14 U3515 ( .A(n3112), .B(n2979), .Z(n2994) );
  HS65_LH_AND2ABX27 U3536 ( .A(n3114), .B(n8573), .Z(n2986) );
  HS65_LL_AOI21X2 U3539 ( .A(n5643), .B(n3888), .C(n3887), .Z(n3889) );
  HS65_LH_OAI21X3 U3544 ( .A(n5201), .B(n5135), .C(n4466), .Z(n4470) );
  HS65_LL_CNBFX21 U3557 ( .A(n5610), .Z(n2859) );
  HS65_LH_IVX9 U3588 ( .A(n9348), .Z(n9349) );
  HS65_LL_NOR2AX3 U3647 ( .A(n3415), .B(n5089), .Z(n4516) );
  HS65_LH_NOR2X6 U3654 ( .A(n2842), .B(n5376), .Z(n4049) );
  HS65_LL_OAI211X8 U3662 ( .A(n7868), .B(n3398), .C(n3397), .D(n3396), .Z(
        n3401) );
  HS65_LH_IVX2 U3721 ( .A(n5127), .Z(n5133) );
  HS65_LH_IVX2 U3736 ( .A(n5474), .Z(n5475) );
  HS65_LH_IVX2 U3779 ( .A(n4050), .Z(n5084) );
  HS65_LH_NAND2X2 U3828 ( .A(n3892), .B(n5295), .Z(n5302) );
  HS65_LH_IVX2 U3877 ( .A(n3967), .Z(n3968) );
  HS65_LH_IVX2 U3924 ( .A(n5299), .Z(n5468) );
  HS65_LH_IVX2 U3958 ( .A(n5186), .Z(n3720) );
  HS65_LH_NAND2X4 U3961 ( .A(n4147), .B(n2848), .Z(n5327) );
  HS65_LH_NAND3X2 U3965 ( .A(n4749), .B(n4870), .C(n4748), .Z(n4760) );
  HS65_LH_NAND3X2 U3966 ( .A(n5563), .B(n5502), .C(n5501), .Z(n5528) );
  HS65_LH_OAI21X2 U4000 ( .A(n5350), .B(n5349), .C(n5348), .Z(n5351) );
  HS65_LH_IVX2 U4042 ( .A(n3665), .Z(n3667) );
  HS65_LH_IVX2 U4099 ( .A(n3836), .Z(n3783) );
  HS65_LH_NAND2X2 U4111 ( .A(n4717), .B(n9342), .Z(n3183) );
  HS65_LH_OR2X4 U4118 ( .A(n4700), .B(n4795), .Z(n3665) );
  HS65_LH_NAND2X2 U4122 ( .A(n5618), .B(n5617), .Z(n5619) );
  HS65_LH_IVX2 U4151 ( .A(n4917), .Z(n3895) );
  HS65_LH_NAND2X2 U4167 ( .A(\sub_x_53/A[23] ), .B(n4351), .Z(n3603) );
  HS65_LH_NAND2X2 U4197 ( .A(n3721), .B(n3720), .Z(n3722) );
  HS65_LH_IVX2 U4203 ( .A(n5346), .Z(n4709) );
  HS65_LH_NOR3X1 U4213 ( .A(n5543), .B(n5542), .C(n5541), .Z(n5561) );
  HS65_LH_CBI4I1X3 U4217 ( .A(n5316), .B(n5315), .C(n5325), .D(n5314), .Z(
        n5485) );
  HS65_LH_IVX2 U4218 ( .A(n4528), .Z(n4196) );
  HS65_LH_NAND2X2 U4221 ( .A(n3494), .B(n3493), .Z(n3495) );
  HS65_LH_NOR2AX3 U4225 ( .A(n3526), .B(n3525), .Z(n3527) );
  HS65_LH_AOI21X2 U4232 ( .A(n5207), .B(n5139), .C(n4853), .Z(n4854) );
  HS65_LH_NAND2X2 U4233 ( .A(n3665), .B(n3594), .Z(n3553) );
  HS65_LH_NAND2X2 U4236 ( .A(n3327), .B(n9177), .Z(n3222) );
  HS65_LH_NAND2X2 U4243 ( .A(n3482), .B(n3939), .Z(n3941) );
  HS65_LHS_XNOR2X3 U4248 ( .A(n8942), .B(\u_DataPath/jaddr_i [21]), .Z(n7108)
         );
  HS65_LH_NOR2X2 U4250 ( .A(n5652), .B(n4582), .Z(n3903) );
  HS65_LH_NOR2X2 U4252 ( .A(n4711), .B(n4582), .Z(n4524) );
  HS65_LH_NOR2X2 U4256 ( .A(n5241), .B(n4185), .Z(n4186) );
  HS65_LH_NAND2X2 U4259 ( .A(\sub_x_53/A[27] ), .B(n4976), .Z(n3684) );
  HS65_LH_AOI21X2 U4264 ( .A(n3368), .B(n4917), .C(n3367), .Z(n3369) );
  HS65_LH_NAND2X2 U4269 ( .A(n4516), .B(n4943), .Z(n4149) );
  HS65_LH_NAND2X2 U4270 ( .A(n9221), .B(n9222), .Z(n4283) );
  HS65_LH_OAI21X2 U4288 ( .A(n4320), .B(n4319), .C(n4318), .Z(n4321) );
  HS65_LH_OAI21X2 U4304 ( .A(n4066), .B(n4490), .C(n6123), .Z(n4072) );
  HS65_LH_AOI21X2 U4311 ( .A(n6123), .B(n4806), .C(n4460), .Z(n4461) );
  HS65_LH_IVX2 U4345 ( .A(n4381), .Z(n4383) );
  HS65_LH_IVX2 U4348 ( .A(n5260), .Z(n4251) );
  HS65_LL_NAND3X2 U4354 ( .A(n5246), .B(n5245), .C(n5244), .Z(n5247) );
  HS65_LH_NAND2AX4 U4366 ( .A(n3456), .B(n3455), .Z(n3458) );
  HS65_LH_IVX2 U4392 ( .A(n5603), .Z(n5604) );
  HS65_LH_OAI21X2 U4434 ( .A(n5789), .B(n5786), .C(n5788), .Z(n5761) );
  HS65_LH_NAND2X2 U4454 ( .A(n3474), .B(n4588), .Z(n3959) );
  HS65_LH_NAND3X2 U4492 ( .A(n7108), .B(n7107), .C(n7106), .Z(n7109) );
  HS65_LH_NOR2X2 U4500 ( .A(n5179), .B(n3294), .Z(n4801) );
  HS65_LH_IVX2 U4504 ( .A(n4622), .Z(n4623) );
  HS65_LH_NAND2X2 U4517 ( .A(\lte_x_59/B[15] ), .B(n2864), .Z(n3833) );
  HS65_LH_NAND2X2 U4542 ( .A(n3426), .B(n4491), .Z(n3979) );
  HS65_LH_IVX2 U4545 ( .A(n4742), .Z(n3534) );
  HS65_LH_IVX2 U4559 ( .A(n3979), .Z(n3757) );
  HS65_LL_AOI12X2 U4573 ( .A(n4708), .B(n4707), .C(n4706), .Z(n4736) );
  HS65_LH_NOR2X2 U4576 ( .A(n3788), .B(n4895), .Z(n3590) );
  HS65_LH_OAI21X2 U4578 ( .A(n6070), .B(n5976), .C(n5978), .Z(n5927) );
  HS65_LH_OAI21X2 U4602 ( .A(n2873), .B(n9346), .C(n4489), .Z(n4493) );
  HS65_LH_IVX2 U4606 ( .A(n4328), .Z(n4329) );
  HS65_LH_NAND2X2 U4607 ( .A(n4873), .B(n4951), .Z(n4065) );
  HS65_LH_NAND2X2 U4611 ( .A(n4383), .B(n4382), .Z(n4387) );
  HS65_LH_NAND2X2 U4625 ( .A(n5272), .B(n5275), .Z(n4248) );
  HS65_LH_NAND2X2 U4633 ( .A(n9285), .B(n8399), .Z(n8291) );
  HS65_LH_NAND2X2 U4638 ( .A(n9175), .B(n9227), .Z(n5884) );
  HS65_LH_AO22X4 U4653 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][0] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][0] ), .Z(n7443)
         );
  HS65_LH_AO22X4 U4701 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][28] ), .B(n7522), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][28] ), .Z(n7503)
         );
  HS65_LH_AOI22X1 U4705 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][5] ), .B(n7286), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][5] ), .D(
        n7285), .Z(n6938) );
  HS65_LH_AO22X4 U4768 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][24] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][24] ), .D(
        n7586), .Z(n7562) );
  HS65_LH_AO22X4 U4820 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][26] ), .B(n7522), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][26] ), .Z(n7328)
         );
  HS65_LH_AO22X4 U4832 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][3] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][3] ), .Z(n7401)
         );
  HS65_LH_NOR2X2 U4842 ( .A(n7658), .B(n7657), .Z(n7684) );
  HS65_LH_AOI22X1 U4846 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][30] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][30] ), .D(
        n2888), .Z(n6129) );
  HS65_LH_IVX2 U4848 ( .A(n5824), .Z(n5825) );
  HS65_LH_OAI22X1 U4855 ( .A(n7112), .B(n7111), .C(n7110), .D(n7109), .Z(n7113) );
  HS65_LH_AOI22X1 U4864 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][2] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][2] ), .D(n2889), .Z(n6960) );
  HS65_LH_AOI22X1 U4868 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][21] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][21] ), .D(
        n2889), .Z(n7590) );
  HS65_LH_AO22X4 U4870 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[7][16] ), .B(n7587), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[12][16] ), .D(
        n7586), .Z(n7542) );
  HS65_LH_AO22X4 U4877 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][29] ), .B(n7522), 
        .C(n6752), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][29] ), .Z(n7529)
         );
  HS65_LH_AO22X4 U4880 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][20] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][20] ), .Z(n7483)
         );
  HS65_LH_AOI22X1 U4889 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][30] ), .B(n7580), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][30] ), .D(
        n7579), .Z(n7417) );
  HS65_LH_AO22X4 U4894 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[31][14] ), .B(n7602), 
        .C(n7601), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][14] ), .Z(n7381)
         );
  HS65_LH_AOI22X1 U4895 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][14] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][14] ), .D(
        n2891), .Z(n7370) );
  HS65_LH_AOI22X1 U4896 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[14][4] ), .B(n7415), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[10][4] ), .D(
        n2891), .Z(n7350) );
  HS65_LH_NOR2X6 U4897 ( .A(n6350), .B(n6352), .Z(n6966) );
  HS65_LH_NOR2X9 U4898 ( .A(n6148), .B(n6152), .Z(n6426) );
  HS65_LH_BFX4 U4902 ( .A(n6637), .Z(n7284) );
  HS65_LH_AO22X4 U4905 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][2] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][2] ), .D(n6619), .Z(n6555) );
  HS65_LH_AOI22X1 U4915 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][25] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][25] ), .D(
        n6625), .Z(n7149) );
  HS65_LH_AO22X4 U4921 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[27][9] ), .B(n7277), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[25][9] ), .D(
        n6629), .Z(n7127) );
  HS65_LH_AO22X4 U4923 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[4][28] ), .B(n7293), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[13][28] ), .D(
        n7292), .Z(n6921) );
  HS65_LH_AOI22X1 U4933 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][17] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][17] ), .D(
        n7294), .Z(n6900) );
  HS65_LH_AOI22X1 U4934 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][31] ), .D(
        n6384), .Z(n6880) );
  HS65_LH_AOI22X1 U4944 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][31] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][31] ), .D(
        n7264), .Z(n6870) );
  HS65_LH_AOI22X1 U4945 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[15][18] ), .B(n7265), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[11][18] ), .D(
        n2888), .Z(n6652) );
  HS65_LH_AO22X4 U4949 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[10][20] ), .B(n6927), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[5][20] ), .D(
        n7266), .Z(n6848) );
  HS65_LH_AO22X4 U4951 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][29] ), .B(n9375), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][29] ), .D(
        n7267), .Z(n7268) );
  HS65_LH_AOI22X1 U4957 ( .A(n3426), .B(n4886), .C(n4836), .D(n4873), .Z(n3556) );
  HS65_LH_AOI22X1 U4969 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][8] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ), .D(n7516), 
        .Z(n6774) );
  HS65_LH_AOI22X1 U5038 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][11] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][11] ), .D(
        n6625), .Z(n6251) );
  HS65_LH_AO22X4 U5042 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][31] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][31] ), .D(
        n7318), .Z(n6677) );
  HS65_LH_AO22X4 U5108 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][6] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][6] ), .Z(n7255)
         );
  HS65_LH_AO22X4 U5120 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][21] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][21] ), .D(
        n6637), .Z(n6195) );
  HS65_LH_AO22X4 U5137 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][17] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][17] ), .Z(n6818)
         );
  HS65_LH_AO22X4 U5149 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][16] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][16] ), .D(
        n6637), .Z(n6175) );
  HS65_LH_AOI22X1 U5207 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[21][23] ), .B(n7524), 
        .C(n7593), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[20][23] ), .Z(n7233)
         );
  HS65_LH_AOI22X1 U5208 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][1] ), .B(n7585), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[1][1] ), .D(n2889), .Z(n6833) );
  HS65_LH_AOI22X1 U5237 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][27] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][27] ), .D(
        n6625), .Z(n6211) );
  HS65_LH_AO22X4 U5270 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[11][19] ), .B(n7578), 
        .C(n7310), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[5][19] ), .Z(n6742)
         );
  HS65_LH_AO22X4 U5293 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][18] ), .B(n7580), 
        .C(n7579), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[2][18] ), .Z(n6327)
         );
  HS65_LH_AOI22X1 U5344 ( .A(n7434), .B(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[13][7] ), .C(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[6][7] ), .D(n7516), 
        .Z(n6726) );
  HS65_LH_AOI22X1 U5355 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][22] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][22] ), .D(
        n6625), .Z(n6271) );
  HS65_LH_AOI22X1 U5395 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[26][24] ), .B(n7273), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[29][24] ), .D(
        n6625), .Z(n6291) );
  HS65_LH_AO22X4 U5453 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][5] ), .B(n7517), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[4][5] ), .D(n7318), .Z(n6704) );
  HS65_LH_AO22X4 U5473 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][12] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][12] ), .Z(n6798)
         );
  HS65_LH_AO22X4 U5496 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ), .B(n7170), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[23][13] ), .D(
        n6637), .Z(n7174) );
  HS65_LH_AOI22X1 U5531 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][14] ), .B(n6376), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[21][14] ), .D(
        n7285), .Z(n6314) );
  HS65_LH_AOI22X1 U5578 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][19] ), .D(
        n7171), .Z(n6523) );
  HS65_LH_AO22X4 U5632 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][7] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][7] ), .D(n7291), .Z(n6450) );
  HS65_LH_AO22X4 U5638 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][12] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][12] ), .D(
        n7291), .Z(n6550) );
  HS65_LH_AOI22X1 U5639 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][6] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][6] ), .D(n7294), .Z(n6488) );
  HS65_LH_AOI22X1 U5650 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[8][3] ), .B(n7297), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[0][3] ), .D(n6942), .Z(n6587) );
  HS65_LH_AOI22X1 U5651 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][3] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][3] ), .D(
        n7264), .Z(n6578) );
  HS65_LH_AOI22X1 U5652 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[12][26] ), .B(n6595), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[14][26] ), .D(
        n7264), .Z(n6498) );
  HS65_LH_AO22X4 U5657 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][8] ), .B(n9374), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[6][8] ), .D(n7267), .Z(n6455) );
  HS65_LH_AOI22X1 U5672 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[24][1] ), .B(n6370), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[28][1] ), .D(
        n6600), .Z(n6604) );
  HS65_LH_AO22X4 U5684 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[9][9] ), .B(n7580), 
        .C(n7579), .D(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][9] ), .Z(n7016) );
  HS65_LH_AOI22X1 U5708 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[16][22] ), .B(n6754), 
        .C(n7594), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[22][22] ), .Z(n7004)
         );
  HS65_LH_AO22X4 U5709 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][4] ), .B(n6426), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][4] ), .D(n7291), .Z(n6645) );
  HS65_LH_IVX2 U5710 ( .A(n3747), .Z(n3748) );
  HS65_LH_NAND2X2 U5711 ( .A(n5131), .B(n4937), .Z(n4959) );
  HS65_LH_NAND2X2 U5723 ( .A(n9183), .B(n9232), .Z(n5777) );
  HS65_LH_NAND2X2 U5725 ( .A(n9342), .B(n9218), .Z(n5797) );
  HS65_LH_OR2X4 U5744 ( .A(n9342), .B(n9210), .Z(n5910) );
  HS65_LH_NAND2X2 U5746 ( .A(n9224), .B(n9226), .Z(n5687) );
  HS65_LH_NOR2X2 U5751 ( .A(n9030), .B(n9223), .Z(n5836) );
  HS65_LH_NOR2AX3 U5755 ( .A(n4299), .B(n4298), .Z(n4300) );
  HS65_LH_OA112X4 U5764 ( .A(n9248), .B(n8880), .C(n8400), .D(n9086), .Z(n9382) );
  HS65_LH_IVX2 U5786 ( .A(n4073), .Z(n4074) );
  HS65_LH_NAND2X2 U5796 ( .A(n5131), .B(n4868), .Z(n4869) );
  HS65_LH_OA12X4 U5801 ( .A(n9122), .B(n8453), .C(n7913), .Z(n9390) );
  HS65_LH_IVX2 U5803 ( .A(n5832), .Z(n5892) );
  HS65_LH_NAND2X2 U5807 ( .A(n5884), .B(n5883), .Z(n5889) );
  HS65_LH_NAND2X2 U5821 ( .A(n4187), .B(n3407), .Z(n3408) );
  HS65_LH_NAND2X2 U5842 ( .A(n4573), .B(n4539), .Z(n4540) );
  HS65_LH_NAND3X2 U5849 ( .A(n2977), .B(n2978), .C(n2976), .Z(n2985) );
  HS65_LH_NAND2X2 U5918 ( .A(n2896), .B(n3226), .Z(n6124) );
  HS65_LH_IVX2 U5926 ( .A(\u_DataPath/dataOut_exe_i [12]), .Z(n3256) );
  HS65_LH_AO22X4 U5945 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][15] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][15] ), .Z(n7195)
         );
  HS65_LH_AO22X4 U5962 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[19][10] ), .B(n7522), 
        .C(n7439), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[23][10] ), .Z(n7215)
         );
  HS65_LH_AOI22X1 U5977 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ), .B(n2887), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[22][0] ), .D(
        n7171), .Z(n6422) );
  HS65_LH_AO22X4 U5999 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[1][10] ), .B(n2884), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[2][10] ), .D(
        n7291), .Z(n6409) );
  HS65_LH_AOI22X1 U6004 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[3][15] ), .B(n6941), 
        .C(\u_DataPath/u_decode_unit/reg_file0/bank_register[7][15] ), .D(
        n7294), .Z(n6387) );
  HS65_LH_OR4X4 U6007 ( .A(n7152), .B(n7151), .C(n2882), .D(n2883), .Z(n7158)
         );
  HS65_LH_NAND2X2 U6023 ( .A(n5643), .B(n4826), .Z(n4827) );
  HS65_LH_OAI21X2 U6028 ( .A(n4803), .B(n4954), .C(n4802), .Z(n4814) );
  HS65_LH_AOI22X1 U6038 ( .A(n5131), .B(n4617), .C(n4887), .D(n4616), .Z(n4618) );
  HS65_LH_IVX2 U6057 ( .A(n7693), .Z(n7738) );
  HS65_LH_IVX2 U6130 ( .A(n8122), .Z(n7761) );
  HS65_LH_NAND2X2 U6133 ( .A(n5624), .B(n4816), .Z(n3568) );
  HS65_LH_IVX2 U6148 ( .A(n7688), .Z(n7771) );
  HS65_LL_OAI112X3 U6151 ( .A(n2920), .B(n5596), .C(n5595), .D(n5594), .Z(
        n5712) );
  HS65_LH_NAND2X2 U6173 ( .A(n4331), .B(n3130), .Z(n3393) );
  HS65_LH_IVX2 U6222 ( .A(\u_DataPath/dataOut_exe_i [28]), .Z(n3127) );
  HS65_LH_NAND2X2 U6228 ( .A(n5877), .B(n6031), .Z(n5830) );
  HS65_LH_AOI21X2 U6239 ( .A(n5866), .B(n5868), .C(n5821), .Z(n5822) );
  HS65_LH_NAND2X2 U6256 ( .A(n8911), .B(n9202), .Z(n5920) );
  HS65_LH_NAND2X2 U6273 ( .A(n9145), .B(n9224), .Z(n5959) );
  HS65_LH_OAI21X2 U6295 ( .A(n5995), .B(n6000), .C(n5997), .Z(n6015) );
  HS65_LH_IVX2 U6318 ( .A(n6019), .Z(n6020) );
  HS65_LH_NAND2X2 U6319 ( .A(n8967), .B(n9220), .Z(n6064) );
  HS65_LH_NOR2X2 U6327 ( .A(n9177), .B(n9229), .Z(n6078) );
  HS65_LH_OR2X4 U6351 ( .A(n8911), .B(n9205), .Z(n6117) );
  HS65_LH_IVX2 U6354 ( .A(n7728), .Z(n7730) );
  HS65_LH_NAND2X2 U6368 ( .A(n7631), .B(n4249), .Z(n4282) );
  HS65_LH_OAI21X2 U6385 ( .A(n5173), .B(n5172), .C(n5171), .Z(n5191) );
  HS65_LH_NAND2X2 U6415 ( .A(n5688), .B(n7729), .Z(n7720) );
  HS65_LH_NAND3X2 U6419 ( .A(Data_out_fromRAM[31]), .B(n8270), .C(n8576), .Z(
        n7346) );
  HS65_LH_OR2X4 U6445 ( .A(n8332), .B(n3340), .Z(n3081) );
  HS65_LH_NOR2X2 U6446 ( .A(n8799), .B(n3403), .Z(n3100) );
  HS65_LH_NAND2X2 U6458 ( .A(n9365), .B(n9040), .Z(n8413) );
  HS65_LH_AOI22X1 U6506 ( .A(n8868), .B(n9144), .C(n9368), .D(n9000), .Z(n8419) );
  HS65_LH_IVX2 U6541 ( .A(n2985), .Z(n2979) );
  HS65_LH_NAND2X2 U6543 ( .A(n7654), .B(n7749), .Z(n7752) );
  HS65_LH_AO22X4 U6584 ( .A(n9256), .B(n9188), .C(n9133), .D(n8933), .Z(
        \u_DataPath/jump_address_i [22]) );
  HS65_LH_AO22X4 U6607 ( .A(n9053), .B(n9188), .C(n9133), .D(n9080), .Z(
        \u_DataPath/jump_address_i [3]) );
  HS65_LH_AO22X4 U6686 ( .A(n8937), .B(n9109), .C(n9188), .D(n9092), .Z(
        \u_DataPath/jump_address_i [0]) );
  HS65_LH_IVX2 U6725 ( .A(n7734), .Z(n7778) );
  HS65_LH_IVX2 U6727 ( .A(n6124), .Z(n8504) );
  HS65_LH_NAND2AX4 U6729 ( .A(n8864), .B(n3291), .Z(n8511) );
  HS65_LH_IVX2 U6732 ( .A(n7775), .Z(n8116) );
  HS65_LL_NAND3X2 U6735 ( .A(n4505), .B(n4511), .C(n4510), .Z(n5250) );
  HS65_LH_NOR4ABX2 U6744 ( .A(n6698), .B(n6697), .C(n6696), .D(n6695), .Z(
        n8158) );
  HS65_LH_NOR4ABX2 U6746 ( .A(n6738), .B(n6737), .C(n6736), .D(n6735), .Z(
        n8180) );
  HS65_LH_NAND2X2 U6749 ( .A(n7631), .B(n4649), .Z(n4650) );
  HS65_LHS_XNOR2X3 U6757 ( .A(n3952), .B(n3951), .Z(n4000) );
  HS65_LH_NAND2X4 U6763 ( .A(n5712), .B(n5711), .Z(n5715) );
  HS65_LH_NAND2X2 U6793 ( .A(n6047), .B(n6046), .Z(n6048) );
  HS65_LH_IVX2 U6831 ( .A(n6051), .Z(n6101) );
  HS65_LH_NAND2X2 U6837 ( .A(n5989), .B(n5787), .Z(n5994) );
  HS65_LH_NOR2X2 U6866 ( .A(n7753), .B(n7752), .Z(n7655) );
  HS65_LH_NOR2X2 U6869 ( .A(n7686), .B(n7755), .Z(n7687) );
  HS65_LH_OAI21X2 U6886 ( .A(n6090), .B(n6089), .C(n6088), .Z(n6091) );
  HS65_LH_IVX2 U6892 ( .A(n9223), .Z(n7791) );
  HS65_LH_NAND3X2 U6907 ( .A(opcode_i[1]), .B(n7643), .C(n7642), .Z(n8047) );
  HS65_LH_NAND2X2 U6908 ( .A(n4485), .B(n4484), .Z(n4486) );
  HS65_LH_NOR3X1 U6956 ( .A(n5191), .B(n5190), .C(n5189), .Z(n5225) );
  HS65_LH_NOR2X2 U6958 ( .A(n8850), .B(n3403), .Z(n3250) );
  HS65_LH_OAI21X2 U6967 ( .A(n7775), .B(n7683), .C(n7682), .Z(n7740) );
  HS65_LH_IVX2 U7003 ( .A(n8236), .Z(n7117) );
  HS65_LHS_XOR2X3 U7022 ( .A(n7785), .B(n7784), .Z(\u_DataPath/pc_4_i [30]) );
  HS65_LH_AO22X4 U7028 ( .A(n9192), .B(n8862), .C(n8690), .D(n9240), .Z(
        \u_DataPath/pc4_to_idexreg_i [0]) );
  HS65_LHS_XOR2X3 U7038 ( .A(n2829), .B(n7747), .Z(\u_DataPath/pc_4_i [9]) );
  HS65_LH_IVX2 U7050 ( .A(Data_out_fromRAM[28]), .Z(n8417) );
  HS65_LH_AO22X4 U7052 ( .A(n9254), .B(n8807), .C(n9240), .D(n8963), .Z(
        \u_DataPath/pc4_to_idexreg_i [6]) );
  HS65_LH_AO22X4 U7090 ( .A(n8782), .B(n9253), .C(n9312), .D(n9142), .Z(
        \u_DataPath/immediate_ext_dec_i [9]) );
  HS65_LH_NOR4ABX2 U7112 ( .A(n7223), .B(n7222), .C(n7221), .D(n7220), .Z(
        n8181) );
  HS65_LH_AO22X4 U7141 ( .A(n8770), .B(n9252), .C(n9305), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [2]) );
  HS65_LH_AO22X4 U7150 ( .A(n8774), .B(n9252), .C(n9304), .D(n9069), .Z(
        \u_DataPath/immediate_ext_dec_i [1]) );
  HS65_LHS_XNOR2X3 U7157 ( .A(n2833), .B(n7749), .Z(\u_DataPath/pc_4_i [10])
         );
  HS65_LHS_XOR2X3 U7202 ( .A(n2823), .B(n7750), .Z(\u_DataPath/pc_4_i [11]) );
  HS65_LHS_XNOR2X3 U7243 ( .A(n6120), .B(n6119), .Z(
        \u_DataPath/u_execute/resAdd1_i [28]) );
  HS65_LHS_XNOR2X3 U7244 ( .A(n7717), .B(n7716), .Z(
        \u_DataPath/u_execute/link_value_i [17]) );
  HS65_LHS_XOR2X3 U7291 ( .A(n7791), .B(n7790), .Z(
        \u_DataPath/u_execute/link_value_i [5]) );
  HS65_LH_IVX2 U7296 ( .A(n8298), .Z(n8299) );
  HS65_LH_IVX2 U7322 ( .A(n8576), .Z(n8271) );
  HS65_LH_IVX2 U7332 ( .A(n3109), .Z(n8578) );
  HS65_LH_IVX2 U7342 ( .A(Data_out_fromRAM[23]), .Z(n8360) );
  HS65_LH_IVX18 U7385 ( .A(n2842), .Z(n4675) );
  HS65_LH_NAND2X7 U7398 ( .A(n5626), .B(n5625), .Z(n5640) );
  HS65_LL_NAND3X6 U7412 ( .A(n8476), .B(n8477), .C(n2918), .Z(n5163) );
  HS65_LH_NAND2AX4 U7429 ( .A(n3282), .B(n3368), .Z(n3370) );
  HS65_LL_AND2X4 U7445 ( .A(n8473), .B(n8472), .Z(n2918) );
  HS65_LL_NOR2AX6 U7464 ( .A(n3948), .B(n3947), .Z(n8473) );
  HS65_LL_NAND2AX7 U7476 ( .A(n2921), .B(n3235), .Z(n4683) );
  HS65_LL_OAI21X2 U7478 ( .A(n4427), .B(n2859), .C(n4426), .Z(n4428) );
  HS65_LL_CNBFX17 U7534 ( .A(\u_DataPath/cw_towb_i [0]), .Z(n3404) );
  HS65_LH_IVX9 U7558 ( .A(n9431), .Z(n3285) );
  HS65_LL_NAND2X7 U7568 ( .A(n7874), .B(n5683), .Z(n5684) );
  HS65_LL_NOR2X9 U7580 ( .A(n5678), .B(n5677), .Z(n7853) );
  HS65_LL_NOR2X6 U7601 ( .A(n4793), .B(n4792), .Z(n4832) );
  HS65_LHS_XOR2X3 U7616 ( .A(n4562), .B(n2897), .Z(n4563) );
  HS65_LL_NAND2X4 U7623 ( .A(n5597), .B(n5712), .Z(n5600) );
  HS65_LL_NAND3X6 U7644 ( .A(n8461), .B(n8459), .C(n5283), .Z(n5601) );
  HS65_LL_BFX9 U7675 ( .A(n9066), .Z(n9347) );
  HS65_LL_NAND2AX21 U7712 ( .A(n5163), .B(n5162), .Z(n5683) );
  HS65_LHS_XOR2X3 U7717 ( .A(n3101), .B(n4997), .Z(n4774) );
  HS65_LL_AOI21X6 U7756 ( .A(n5285), .B(n3697), .C(n3696), .Z(n8461) );
  HS65_LH_AO22X4 U7760 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][15] ), .B(n7523), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][15] ), .Z(n7194)
         );
  HS65_LH_AO22X4 U7784 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][8] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][8] ), .Z(n6777)
         );
  HS65_LH_AO22X4 U7814 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][23] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][23] ), .Z(n7234)
         );
  HS65_LH_AO22X4 U7816 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][6] ), .B(n7523), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][6] ), .Z(n7254)
         );
  HS65_LH_AO22X4 U7819 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][31] ), .B(n7523), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][31] ), .Z(n6687)
         );
  HS65_LH_AO22X4 U7830 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][7] ), .B(n7523), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][7] ), .Z(n6729)
         );
  HS65_LH_AO22X4 U7846 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][30] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][30] ), .Z(n7422)
         );
  HS65_LH_AO22X4 U7868 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][20] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][20] ), .Z(n7482)
         );
  HS65_LH_AO22X4 U7871 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][3] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][3] ), .Z(n7397)
         );
  HS65_LH_AO22X4 U7881 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][28] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][28] ), .Z(n7502)
         );
  HS65_LH_AO22X4 U7900 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][14] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][14] ), .Z(n7377)
         );
  HS65_LH_AO22X4 U7901 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][29] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][29] ), .Z(n7528)
         );
  HS65_LH_AO22X4 U7902 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][0] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][0] ), .Z(n7442)
         );
  HS65_LH_AO22X4 U7903 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][13] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][13] ), .Z(n6986)
         );
  HS65_LH_AO22X4 U7904 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][22] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][22] ), .Z(n7006)
         );
  HS65_LH_AO22X4 U8092 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][9] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][9] ), .Z(n7026)
         );
  HS65_LH_AO22X4 U8133 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][11] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][11] ), .Z(n7066)
         );
  HS65_LH_AO22X4 U8136 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][25] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][25] ), .Z(n7046)
         );
  HS65_LH_AO22X4 U8152 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][19] ), .B(n6681), 
        .C(n7592), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][19] ), .Z(n6757)
         );
  HS65_LH_AO22X4 U8162 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][18] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][18] ), .Z(n6345)
         );
  HS65_LH_AO22X4 U8169 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][12] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][12] ), .Z(n6797)
         );
  HS65_LH_AO22X4 U8175 ( .A(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[17][1] ), .B(n7523), 
        .C(n6682), .D(
        \u_DataPath/u_decode_unit/reg_file0/bank_register[18][1] ), .Z(n6837)
         );
  HS65_LHS_XNOR2X3 U8179 ( .A(n4598), .B(n4597), .Z(n4599) );
  HS65_LL_AND2X9 U8184 ( .A(n3397), .B(n3293), .Z(n4805) );
  HS65_LL_NOR2X5 U8198 ( .A(n5161), .B(n5710), .Z(n5162) );
  HS65_LL_NAND3AX6 U8203 ( .A(n5686), .B(n8474), .C(n8475), .Z(n5161) );
  HS65_LL_NOR3X4 U8219 ( .A(n7867), .B(n4302), .C(n5708), .Z(n4456) );
  HS65_LH_NAND2X7 U8277 ( .A(\lte_x_59/B[8] ), .B(n4551), .Z(n3867) );
  HS65_LH_AOI12X2 U8297 ( .A(n3688), .B(n5211), .C(n3687), .Z(n3689) );
  HS65_LL_CNIVX7 U8319 ( .A(n4427), .Z(n2867) );
  HS65_LH_IVX4 U8332 ( .A(n9348), .Z(n9352) );
  HS65_LH_IVX7 U8339 ( .A(n9376), .Z(n4717) );
  HS65_LH_CNIVX3 U8349 ( .A(\u_DataPath/jaddr_i [20]), .Z(n2881) );
  HS65_LH_NOR2X5 U8351 ( .A(n5054), .B(n5053), .Z(n5299) );
  HS65_LL_NAND3X2 U8361 ( .A(n3871), .B(n3870), .C(n3869), .Z(n5143) );
endmodule

