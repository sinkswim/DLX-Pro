
module mmu_out_dram ( data_ram, mem_op, nibble, unaligned, data_read );
  input [31:0] data_ram;
  input [5:0] mem_op;
  input [1:0] nibble;
  output [31:0] data_read;
  input unaligned;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n3, n4;

  NAND3_X1 U100 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n42) );
  NAND3_X1 U102 ( .A1(n101), .A2(n100), .A3(n102), .ZN(n46) );
  XOR2_X1 U103 ( .A(mem_op[3]), .B(mem_op[0]), .Z(n102) );
  NOR4_X1 U2 ( .A1(n101), .A2(mem_op[0]), .A3(mem_op[2]), .A4(mem_op[3]), .ZN(
        n93) );
  OR2_X1 U3 ( .A1(n49), .A2(n92), .ZN(n35) );
  INV_X1 U4 ( .A(n91), .ZN(n96) );
  OR2_X1 U5 ( .A1(n86), .A2(nibble[0]), .ZN(n88) );
  OAI22_X1 U6 ( .A1(n96), .A2(n97), .B1(n46), .B2(n98), .ZN(n53) );
  INV_X1 U7 ( .A(n93), .ZN(n97) );
  NAND2_X1 U8 ( .A1(nibble[0]), .A2(n86), .ZN(n98) );
  NAND2_X1 U9 ( .A1(n78), .A2(n43), .ZN(n61) );
  OAI21_X1 U10 ( .B1(n46), .B2(n99), .A(n92), .ZN(n52) );
  NAND2_X1 U11 ( .A1(nibble[1]), .A2(nibble[0]), .ZN(n99) );
  NOR2_X1 U12 ( .A1(n46), .A2(n88), .ZN(n50) );
  NOR2_X1 U13 ( .A1(n46), .A2(n96), .ZN(n51) );
  NAND3_X1 U14 ( .A1(n43), .A2(n91), .A3(n93), .ZN(n33) );
  INV_X1 U15 ( .A(n43), .ZN(n49) );
  NOR2_X1 U16 ( .A1(nibble[0]), .A2(nibble[1]), .ZN(n91) );
  BUF_X1 U17 ( .A(n37), .Z(n3) );
  BUF_X1 U18 ( .A(n37), .Z(n4) );
  AOI21_X1 U19 ( .B1(n96), .B2(n93), .A(n78), .ZN(n92) );
  INV_X1 U20 ( .A(nibble[1]), .ZN(n86) );
  INV_X1 U21 ( .A(n46), .ZN(n45) );
  OAI221_X1 U22 ( .B1(n60), .B2(n33), .C1(n79), .C2(n35), .A(n3), .ZN(
        data_read[15]) );
  OAI21_X1 U23 ( .B1(n61), .B2(n68), .A(n4), .ZN(data_read[26]) );
  OAI21_X1 U24 ( .B1(n40), .B2(n61), .A(n4), .ZN(data_read[23]) );
  OAI21_X1 U25 ( .B1(n38), .B2(n61), .A(n4), .ZN(data_read[24]) );
  OAI21_X1 U26 ( .B1(n34), .B2(n61), .A(n4), .ZN(data_read[25]) );
  OAI21_X1 U27 ( .B1(n67), .B2(n61), .A(n4), .ZN(data_read[27]) );
  OAI21_X1 U28 ( .B1(n66), .B2(n61), .A(n4), .ZN(data_read[28]) );
  OAI21_X1 U29 ( .B1(n65), .B2(n61), .A(n4), .ZN(data_read[29]) );
  OAI21_X1 U30 ( .B1(n62), .B2(n61), .A(n4), .ZN(data_read[30]) );
  OAI21_X1 U31 ( .B1(n60), .B2(n61), .A(n3), .ZN(data_read[31]) );
  NOR3_X1 U32 ( .A1(unaligned), .A2(mem_op[5]), .A3(mem_op[4]), .ZN(n43) );
  NOR4_X1 U33 ( .A1(n100), .A2(mem_op[0]), .A3(mem_op[1]), .A4(mem_op[3]), 
        .ZN(n78) );
  OAI221_X1 U34 ( .B1(n86), .B2(n87), .C1(n88), .C2(n79), .A(n89), .ZN(n44) );
  NAND2_X1 U35 ( .A1(data_ram[7]), .A2(nibble[0]), .ZN(n87) );
  AOI22_X1 U36 ( .A1(n90), .A2(nibble[0]), .B1(data_ram[31]), .B2(n91), .ZN(
        n89) );
  NOR2_X1 U37 ( .A1(nibble[1]), .A2(n40), .ZN(n90) );
  NAND4_X1 U38 ( .A1(n43), .A2(n44), .A3(mem_op[0]), .A4(n85), .ZN(n37) );
  NOR3_X1 U39 ( .A1(mem_op[1]), .A2(mem_op[3]), .A3(mem_op[2]), .ZN(n85) );
  INV_X1 U40 ( .A(data_ram[23]), .ZN(n40) );
  INV_X1 U41 ( .A(mem_op[2]), .ZN(n100) );
  INV_X1 U42 ( .A(mem_op[1]), .ZN(n101) );
  INV_X1 U43 ( .A(data_ram[31]), .ZN(n60) );
  INV_X1 U44 ( .A(data_ram[26]), .ZN(n68) );
  INV_X1 U45 ( .A(data_ram[15]), .ZN(n79) );
  INV_X1 U46 ( .A(data_ram[24]), .ZN(n38) );
  INV_X1 U47 ( .A(data_ram[25]), .ZN(n34) );
  INV_X1 U48 ( .A(data_ram[27]), .ZN(n67) );
  INV_X1 U49 ( .A(data_ram[28]), .ZN(n66) );
  INV_X1 U50 ( .A(data_ram[29]), .ZN(n65) );
  INV_X1 U51 ( .A(data_ram[30]), .ZN(n62) );
  OAI221_X1 U52 ( .B1(n33), .B2(n38), .C1(n35), .C2(n39), .A(n3), .ZN(
        data_read[8]) );
  INV_X1 U53 ( .A(data_ram[8]), .ZN(n39) );
  OAI221_X1 U54 ( .B1(n33), .B2(n34), .C1(n35), .C2(n36), .A(n3), .ZN(
        data_read[9]) );
  INV_X1 U55 ( .A(data_ram[9]), .ZN(n36) );
  OAI221_X1 U56 ( .B1(n33), .B2(n68), .C1(n35), .C2(n84), .A(n3), .ZN(
        data_read[10]) );
  INV_X1 U57 ( .A(data_ram[10]), .ZN(n84) );
  OAI221_X1 U58 ( .B1(n33), .B2(n67), .C1(n35), .C2(n83), .A(n3), .ZN(
        data_read[11]) );
  INV_X1 U59 ( .A(data_ram[11]), .ZN(n83) );
  OAI221_X1 U60 ( .B1(n33), .B2(n66), .C1(n35), .C2(n82), .A(n3), .ZN(
        data_read[12]) );
  INV_X1 U61 ( .A(data_ram[12]), .ZN(n82) );
  OAI221_X1 U62 ( .B1(n33), .B2(n65), .C1(n35), .C2(n81), .A(n3), .ZN(
        data_read[13]) );
  INV_X1 U63 ( .A(data_ram[13]), .ZN(n81) );
  OAI221_X1 U64 ( .B1(n33), .B2(n62), .C1(n35), .C2(n80), .A(n3), .ZN(
        data_read[14]) );
  INV_X1 U65 ( .A(data_ram[14]), .ZN(n80) );
  OAI221_X1 U66 ( .B1(n40), .B2(n33), .C1(n41), .C2(n35), .A(n42), .ZN(
        data_read[7]) );
  INV_X1 U67 ( .A(data_ram[7]), .ZN(n41) );
  OAI21_X1 U68 ( .B1(n61), .B2(n77), .A(n3), .ZN(data_read[16]) );
  INV_X1 U69 ( .A(data_ram[16]), .ZN(n77) );
  OAI21_X1 U70 ( .B1(n61), .B2(n76), .A(n3), .ZN(data_read[17]) );
  INV_X1 U71 ( .A(data_ram[17]), .ZN(n76) );
  OAI21_X1 U72 ( .B1(n61), .B2(n75), .A(n3), .ZN(data_read[18]) );
  INV_X1 U73 ( .A(data_ram[18]), .ZN(n75) );
  OAI21_X1 U74 ( .B1(n74), .B2(n61), .A(n4), .ZN(data_read[19]) );
  INV_X1 U75 ( .A(data_ram[19]), .ZN(n74) );
  OAI21_X1 U76 ( .B1(n71), .B2(n61), .A(n4), .ZN(data_read[20]) );
  INV_X1 U77 ( .A(data_ram[20]), .ZN(n71) );
  OAI21_X1 U78 ( .B1(n70), .B2(n61), .A(n4), .ZN(data_read[21]) );
  INV_X1 U79 ( .A(data_ram[21]), .ZN(n70) );
  OAI21_X1 U80 ( .B1(n69), .B2(n61), .A(n4), .ZN(data_read[22]) );
  INV_X1 U81 ( .A(data_ram[22]), .ZN(n69) );
  AOI21_X1 U82 ( .B1(n94), .B2(n95), .A(n49), .ZN(data_read[0]) );
  AOI22_X1 U83 ( .A1(n50), .A2(data_ram[8]), .B1(n51), .B2(data_ram[24]), .ZN(
        n95) );
  AOI22_X1 U84 ( .A1(data_ram[0]), .A2(n52), .B1(data_ram[16]), .B2(n53), .ZN(
        n94) );
  AOI21_X1 U85 ( .B1(n72), .B2(n73), .A(n49), .ZN(data_read[1]) );
  AOI22_X1 U86 ( .A1(n50), .A2(data_ram[9]), .B1(n51), .B2(data_ram[25]), .ZN(
        n73) );
  AOI22_X1 U87 ( .A1(data_ram[1]), .A2(n52), .B1(data_ram[17]), .B2(n53), .ZN(
        n72) );
  AOI21_X1 U88 ( .B1(n63), .B2(n64), .A(n49), .ZN(data_read[2]) );
  AOI22_X1 U89 ( .A1(data_ram[2]), .A2(n52), .B1(data_ram[18]), .B2(n53), .ZN(
        n63) );
  AOI22_X1 U90 ( .A1(data_ram[10]), .A2(n50), .B1(data_ram[26]), .B2(n51), 
        .ZN(n64) );
  AOI21_X1 U91 ( .B1(n58), .B2(n59), .A(n49), .ZN(data_read[3]) );
  AOI22_X1 U92 ( .A1(data_ram[3]), .A2(n52), .B1(data_ram[19]), .B2(n53), .ZN(
        n58) );
  AOI22_X1 U93 ( .A1(data_ram[11]), .A2(n50), .B1(data_ram[27]), .B2(n51), 
        .ZN(n59) );
  AOI21_X1 U94 ( .B1(n56), .B2(n57), .A(n49), .ZN(data_read[4]) );
  AOI22_X1 U95 ( .A1(data_ram[4]), .A2(n52), .B1(data_ram[20]), .B2(n53), .ZN(
        n56) );
  AOI22_X1 U96 ( .A1(data_ram[12]), .A2(n50), .B1(data_ram[28]), .B2(n51), 
        .ZN(n57) );
  AOI21_X1 U97 ( .B1(n54), .B2(n55), .A(n49), .ZN(data_read[5]) );
  AOI22_X1 U98 ( .A1(data_ram[5]), .A2(n52), .B1(data_ram[21]), .B2(n53), .ZN(
        n54) );
  AOI22_X1 U99 ( .A1(data_ram[13]), .A2(n50), .B1(data_ram[29]), .B2(n51), 
        .ZN(n55) );
  AOI21_X1 U101 ( .B1(n47), .B2(n48), .A(n49), .ZN(data_read[6]) );
  AOI22_X1 U104 ( .A1(data_ram[6]), .A2(n52), .B1(data_ram[22]), .B2(n53), 
        .ZN(n47) );
  AOI22_X1 U105 ( .A1(data_ram[14]), .A2(n50), .B1(data_ram[30]), .B2(n51), 
        .ZN(n48) );
endmodule


module mmu_in_dram ( mem_op, aligned_address, data, unaligned, nibble, 
        write_op, read_op, mem_address, mem_data, write_byte );
  input [5:0] mem_op;
  input [31:0] aligned_address;
  input [31:0] data;
  output [1:0] nibble;
  output [31:0] mem_address;
  output [31:0] mem_data;
  output unaligned, write_op, read_op, write_byte;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n7, n8, n9, n33, n34;
  assign mem_address[31] = 1'b0;
  assign mem_address[30] = 1'b0;

  BUF_X1 U3 ( .A(n24), .Z(n8) );
  BUF_X1 U4 ( .A(n24), .Z(n7) );
  BUF_X1 U5 ( .A(n24), .Z(n9) );
  NAND2_X1 U6 ( .A1(n12), .A2(n20), .ZN(n24) );
  NOR2_X1 U7 ( .A1(n20), .A2(n13), .ZN(nibble[0]) );
  AND3_X1 U8 ( .A1(n16), .A2(n23), .A3(n15), .ZN(n20) );
  AND2_X1 U9 ( .A1(n10), .A2(n17), .ZN(n12) );
  AND2_X1 U10 ( .A1(n18), .A2(n22), .ZN(n10) );
  OR2_X1 U11 ( .A1(write_byte), .A2(n21), .ZN(write_op) );
  BUF_X1 U12 ( .A(n21), .Z(n34) );
  BUF_X1 U13 ( .A(n21), .Z(n33) );
  INV_X1 U14 ( .A(n23), .ZN(write_byte) );
  NOR3_X1 U15 ( .A1(mem_op[1]), .A2(mem_op[2]), .A3(mem_op[0]), .ZN(n25) );
  NOR3_X1 U16 ( .A1(mem_op[4]), .A2(mem_op[5]), .A3(mem_op[3]), .ZN(n29) );
  OAI22_X1 U17 ( .A1(n10), .A2(n11), .B1(n12), .B2(n13), .ZN(unaligned) );
  INV_X1 U18 ( .A(aligned_address[1]), .ZN(n11) );
  NAND4_X1 U19 ( .A1(mem_op[1]), .A2(n29), .A3(n32), .A4(n31), .ZN(n17) );
  NAND4_X1 U20 ( .A1(mem_op[0]), .A2(n29), .A3(n30), .A4(n31), .ZN(n16) );
  NAND4_X1 U21 ( .A1(mem_op[3]), .A2(n25), .A3(n26), .A4(n27), .ZN(n15) );
  NAND4_X1 U22 ( .A1(mem_op[2]), .A2(n29), .A3(n32), .A4(n30), .ZN(n18) );
  NAND4_X1 U23 ( .A1(mem_op[4]), .A2(n25), .A3(n28), .A4(n27), .ZN(n22) );
  NAND4_X1 U24 ( .A1(mem_op[5]), .A2(n25), .A3(n28), .A4(n26), .ZN(n23) );
  AND2_X1 U25 ( .A1(n19), .A2(aligned_address[1]), .ZN(nibble[1]) );
  OAI21_X1 U26 ( .B1(n17), .B2(aligned_address[0]), .A(n20), .ZN(n19) );
  INV_X1 U27 ( .A(mem_op[3]), .ZN(n28) );
  INV_X1 U28 ( .A(mem_op[0]), .ZN(n32) );
  INV_X1 U29 ( .A(mem_op[2]), .ZN(n31) );
  INV_X1 U30 ( .A(mem_op[1]), .ZN(n30) );
  INV_X1 U31 ( .A(aligned_address[0]), .ZN(n13) );
  INV_X1 U32 ( .A(mem_op[5]), .ZN(n27) );
  INV_X1 U33 ( .A(mem_op[4]), .ZN(n26) );
  NOR3_X1 U34 ( .A1(aligned_address[0]), .A2(aligned_address[1]), .A3(n22), 
        .ZN(n21) );
  NAND4_X1 U35 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(read_op) );
  OR3_X1 U36 ( .A1(aligned_address[0]), .A2(aligned_address[1]), .A3(n18), 
        .ZN(n14) );
  AND2_X1 U37 ( .A1(data[0]), .A2(write_op), .ZN(mem_data[0]) );
  AND2_X1 U38 ( .A1(data[1]), .A2(write_op), .ZN(mem_data[1]) );
  AND2_X1 U39 ( .A1(data[2]), .A2(write_op), .ZN(mem_data[2]) );
  AND2_X1 U40 ( .A1(data[3]), .A2(write_op), .ZN(mem_data[3]) );
  AND2_X1 U41 ( .A1(data[4]), .A2(write_op), .ZN(mem_data[4]) );
  AND2_X1 U42 ( .A1(data[5]), .A2(write_op), .ZN(mem_data[5]) );
  AND2_X1 U43 ( .A1(data[6]), .A2(write_op), .ZN(mem_data[6]) );
  AND2_X1 U44 ( .A1(data[7]), .A2(write_op), .ZN(mem_data[7]) );
  AND2_X1 U45 ( .A1(data[8]), .A2(n33), .ZN(mem_data[8]) );
  AND2_X1 U46 ( .A1(data[9]), .A2(n33), .ZN(mem_data[9]) );
  AND2_X1 U47 ( .A1(data[10]), .A2(n34), .ZN(mem_data[10]) );
  AND2_X1 U48 ( .A1(data[11]), .A2(n34), .ZN(mem_data[11]) );
  AND2_X1 U49 ( .A1(data[12]), .A2(n34), .ZN(mem_data[12]) );
  AND2_X1 U50 ( .A1(data[13]), .A2(n34), .ZN(mem_data[13]) );
  AND2_X1 U51 ( .A1(data[14]), .A2(n34), .ZN(mem_data[14]) );
  AND2_X1 U52 ( .A1(data[15]), .A2(n34), .ZN(mem_data[15]) );
  AND2_X1 U53 ( .A1(data[16]), .A2(n34), .ZN(mem_data[16]) );
  AND2_X1 U54 ( .A1(data[17]), .A2(n34), .ZN(mem_data[17]) );
  AND2_X1 U55 ( .A1(data[18]), .A2(n34), .ZN(mem_data[18]) );
  AND2_X1 U56 ( .A1(data[19]), .A2(n34), .ZN(mem_data[19]) );
  AND2_X1 U57 ( .A1(data[20]), .A2(n34), .ZN(mem_data[20]) );
  AND2_X1 U58 ( .A1(data[21]), .A2(n34), .ZN(mem_data[21]) );
  AND2_X1 U59 ( .A1(data[22]), .A2(n33), .ZN(mem_data[22]) );
  AND2_X1 U60 ( .A1(data[23]), .A2(n33), .ZN(mem_data[23]) );
  AND2_X1 U61 ( .A1(data[24]), .A2(n33), .ZN(mem_data[24]) );
  AND2_X1 U62 ( .A1(data[25]), .A2(n33), .ZN(mem_data[25]) );
  AND2_X1 U63 ( .A1(data[26]), .A2(n33), .ZN(mem_data[26]) );
  AND2_X1 U64 ( .A1(data[27]), .A2(n33), .ZN(mem_data[27]) );
  AND2_X1 U65 ( .A1(data[28]), .A2(n33), .ZN(mem_data[28]) );
  AND2_X1 U66 ( .A1(data[29]), .A2(n33), .ZN(mem_data[29]) );
  AND2_X1 U67 ( .A1(data[30]), .A2(n33), .ZN(mem_data[30]) );
  AND2_X1 U68 ( .A1(data[31]), .A2(n33), .ZN(mem_data[31]) );
  AND2_X1 U69 ( .A1(aligned_address[3]), .A2(n8), .ZN(mem_address[1]) );
  AND2_X1 U70 ( .A1(aligned_address[4]), .A2(n7), .ZN(mem_address[2]) );
  AND2_X1 U71 ( .A1(aligned_address[5]), .A2(n7), .ZN(mem_address[3]) );
  AND2_X1 U72 ( .A1(aligned_address[6]), .A2(n7), .ZN(mem_address[4]) );
  AND2_X1 U73 ( .A1(aligned_address[7]), .A2(n7), .ZN(mem_address[5]) );
  AND2_X1 U74 ( .A1(aligned_address[8]), .A2(n7), .ZN(mem_address[6]) );
  AND2_X1 U75 ( .A1(aligned_address[9]), .A2(n7), .ZN(mem_address[7]) );
  AND2_X1 U76 ( .A1(aligned_address[10]), .A2(n7), .ZN(mem_address[8]) );
  AND2_X1 U77 ( .A1(aligned_address[11]), .A2(n7), .ZN(mem_address[9]) );
  AND2_X1 U78 ( .A1(aligned_address[17]), .A2(n8), .ZN(mem_address[15]) );
  AND2_X1 U79 ( .A1(aligned_address[18]), .A2(n8), .ZN(mem_address[16]) );
  AND2_X1 U80 ( .A1(aligned_address[19]), .A2(n8), .ZN(mem_address[17]) );
  AND2_X1 U81 ( .A1(aligned_address[20]), .A2(n8), .ZN(mem_address[18]) );
  AND2_X1 U82 ( .A1(aligned_address[21]), .A2(n8), .ZN(mem_address[19]) );
  AND2_X1 U83 ( .A1(aligned_address[22]), .A2(n8), .ZN(mem_address[20]) );
  AND2_X1 U84 ( .A1(aligned_address[23]), .A2(n8), .ZN(mem_address[21]) );
  AND2_X1 U85 ( .A1(aligned_address[24]), .A2(n8), .ZN(mem_address[22]) );
  AND2_X1 U86 ( .A1(aligned_address[25]), .A2(n8), .ZN(mem_address[23]) );
  AND2_X1 U87 ( .A1(aligned_address[26]), .A2(n8), .ZN(mem_address[24]) );
  AND2_X1 U88 ( .A1(aligned_address[27]), .A2(n8), .ZN(mem_address[25]) );
  AND2_X1 U89 ( .A1(aligned_address[28]), .A2(n7), .ZN(mem_address[26]) );
  AND2_X1 U90 ( .A1(aligned_address[29]), .A2(n7), .ZN(mem_address[27]) );
  AND2_X1 U91 ( .A1(aligned_address[30]), .A2(n7), .ZN(mem_address[28]) );
  AND2_X1 U92 ( .A1(aligned_address[31]), .A2(n7), .ZN(mem_address[29]) );
  AND2_X1 U93 ( .A1(aligned_address[2]), .A2(n9), .ZN(mem_address[0]) );
  AND2_X1 U94 ( .A1(aligned_address[12]), .A2(n9), .ZN(mem_address[10]) );
  AND2_X1 U95 ( .A1(aligned_address[13]), .A2(n9), .ZN(mem_address[11]) );
  AND2_X1 U96 ( .A1(aligned_address[14]), .A2(n9), .ZN(mem_address[12]) );
  AND2_X1 U97 ( .A1(aligned_address[15]), .A2(n9), .ZN(mem_address[13]) );
  AND2_X1 U98 ( .A1(aligned_address[16]), .A2(n9), .ZN(mem_address[14]) );
endmodule


module ALU_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199;

  XOR2_X1 U55 ( .A(A[30]), .B(n111), .Z(n7) );
  NAND3_X1 U149 ( .A1(n189), .A2(n99), .A3(n96), .ZN(n185) );
  NAND3_X1 U153 ( .A1(n193), .A2(n194), .A3(n195), .ZN(n189) );
  INV_X1 U1 ( .A(n91), .ZN(n88) );
  INV_X1 U2 ( .A(n77), .ZN(n74) );
  INV_X1 U3 ( .A(n63), .ZN(n60) );
  INV_X1 U4 ( .A(n49), .ZN(n46) );
  INV_X1 U5 ( .A(n35), .ZN(n32) );
  INV_X1 U6 ( .A(n21), .ZN(n18) );
  INV_X1 U7 ( .A(EQ), .ZN(NE) );
  NOR2_X1 U8 ( .A1(GT), .A2(LT), .ZN(EQ) );
  NOR2_X1 U9 ( .A1(n179), .A2(n83), .ZN(n82) );
  NOR2_X1 U10 ( .A1(n167), .A2(n69), .ZN(n68) );
  NOR2_X1 U11 ( .A1(n155), .A2(n55), .ZN(n54) );
  NOR2_X1 U12 ( .A1(n143), .A2(n41), .ZN(n40) );
  NOR2_X1 U13 ( .A1(n131), .A2(n27), .ZN(n26) );
  NOR2_X1 U14 ( .A1(n119), .A2(n13), .ZN(n12) );
  OAI211_X1 U15 ( .C1(n117), .C2(n118), .A(n15), .B(n12), .ZN(n114) );
  NAND2_X1 U16 ( .A1(n122), .A2(n123), .ZN(n118) );
  AOI211_X1 U17 ( .C1(n124), .C2(n125), .A(n21), .B(n126), .ZN(n117) );
  INV_X1 U18 ( .A(n16), .ZN(n122) );
  OAI211_X1 U19 ( .C1(n177), .C2(n178), .A(n85), .B(n82), .ZN(n173) );
  NAND2_X1 U20 ( .A1(n182), .A2(n183), .ZN(n178) );
  AOI211_X1 U21 ( .C1(n184), .C2(n185), .A(n91), .B(n186), .ZN(n177) );
  INV_X1 U22 ( .A(n86), .ZN(n182) );
  OAI211_X1 U23 ( .C1(n165), .C2(n166), .A(n71), .B(n68), .ZN(n161) );
  NAND2_X1 U24 ( .A1(n170), .A2(n171), .ZN(n166) );
  AOI211_X1 U25 ( .C1(n172), .C2(n173), .A(n77), .B(n174), .ZN(n165) );
  INV_X1 U26 ( .A(n72), .ZN(n170) );
  OAI211_X1 U27 ( .C1(n153), .C2(n154), .A(n57), .B(n54), .ZN(n149) );
  NAND2_X1 U28 ( .A1(n158), .A2(n159), .ZN(n154) );
  AOI211_X1 U29 ( .C1(n160), .C2(n161), .A(n63), .B(n162), .ZN(n153) );
  INV_X1 U30 ( .A(n58), .ZN(n158) );
  OAI211_X1 U31 ( .C1(n141), .C2(n142), .A(n43), .B(n40), .ZN(n137) );
  NAND2_X1 U32 ( .A1(n146), .A2(n147), .ZN(n142) );
  AOI211_X1 U33 ( .C1(n148), .C2(n149), .A(n49), .B(n150), .ZN(n141) );
  INV_X1 U34 ( .A(n44), .ZN(n146) );
  OAI211_X1 U35 ( .C1(n129), .C2(n130), .A(n29), .B(n26), .ZN(n125) );
  NAND2_X1 U36 ( .A1(n134), .A2(n135), .ZN(n130) );
  AOI211_X1 U37 ( .C1(n136), .C2(n137), .A(n35), .B(n138), .ZN(n129) );
  INV_X1 U38 ( .A(n30), .ZN(n134) );
  AOI21_X1 U39 ( .B1(n92), .B2(n93), .A(n94), .ZN(n87) );
  AOI21_X1 U40 ( .B1(n95), .B2(n96), .A(n97), .ZN(n92) );
  AOI21_X1 U41 ( .B1(n98), .B2(n99), .A(n100), .ZN(n95) );
  AOI21_X1 U42 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  AOI21_X1 U43 ( .B1(n78), .B2(n79), .A(n80), .ZN(n73) );
  AOI21_X1 U44 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  AOI21_X1 U45 ( .B1(n84), .B2(n85), .A(n86), .ZN(n81) );
  AOI21_X1 U46 ( .B1(n87), .B2(n88), .A(n89), .ZN(n84) );
  AOI21_X1 U47 ( .B1(n64), .B2(n65), .A(n66), .ZN(n59) );
  AOI21_X1 U48 ( .B1(n67), .B2(n68), .A(n69), .ZN(n64) );
  AOI21_X1 U49 ( .B1(n70), .B2(n71), .A(n72), .ZN(n67) );
  AOI21_X1 U50 ( .B1(n73), .B2(n74), .A(n75), .ZN(n70) );
  AOI21_X1 U51 ( .B1(n50), .B2(n51), .A(n52), .ZN(n45) );
  AOI21_X1 U52 ( .B1(n53), .B2(n54), .A(n55), .ZN(n50) );
  AOI21_X1 U53 ( .B1(n56), .B2(n57), .A(n58), .ZN(n53) );
  AOI21_X1 U54 ( .B1(n59), .B2(n60), .A(n61), .ZN(n56) );
  AOI21_X1 U56 ( .B1(n36), .B2(n37), .A(n38), .ZN(n31) );
  AOI21_X1 U57 ( .B1(n39), .B2(n40), .A(n41), .ZN(n36) );
  AOI21_X1 U58 ( .B1(n42), .B2(n43), .A(n44), .ZN(n39) );
  AOI21_X1 U59 ( .B1(n45), .B2(n46), .A(n47), .ZN(n42) );
  AOI21_X1 U60 ( .B1(n22), .B2(n23), .A(n24), .ZN(n17) );
  AOI21_X1 U61 ( .B1(n25), .B2(n26), .A(n27), .ZN(n22) );
  AOI21_X1 U62 ( .B1(n28), .B2(n29), .A(n30), .ZN(n25) );
  AOI21_X1 U63 ( .B1(n31), .B2(n32), .A(n33), .ZN(n28) );
  AOI21_X1 U64 ( .B1(n8), .B2(n9), .A(n10), .ZN(n6) );
  AOI21_X1 U65 ( .B1(n11), .B2(n12), .A(n13), .ZN(n8) );
  AOI21_X1 U66 ( .B1(n14), .B2(n15), .A(n16), .ZN(n11) );
  AOI21_X1 U67 ( .B1(n17), .B2(n18), .A(n19), .ZN(n14) );
  NOR2_X1 U68 ( .A1(n190), .A2(n97), .ZN(n96) );
  NOR2_X1 U69 ( .A1(n190), .A2(n94), .ZN(n184) );
  NOR2_X1 U70 ( .A1(n179), .A2(n80), .ZN(n172) );
  NOR2_X1 U71 ( .A1(n167), .A2(n66), .ZN(n160) );
  NOR2_X1 U72 ( .A1(n155), .A2(n52), .ZN(n148) );
  NOR2_X1 U73 ( .A1(n143), .A2(n38), .ZN(n136) );
  NOR2_X1 U74 ( .A1(n131), .A2(n24), .ZN(n124) );
  NOR2_X1 U75 ( .A1(n119), .A2(n10), .ZN(n113) );
  NAND2_X1 U76 ( .A1(n183), .A2(n90), .ZN(n91) );
  NAND2_X1 U77 ( .A1(n171), .A2(n76), .ZN(n77) );
  NAND2_X1 U78 ( .A1(n159), .A2(n62), .ZN(n63) );
  NAND2_X1 U79 ( .A1(n147), .A2(n48), .ZN(n49) );
  NAND2_X1 U80 ( .A1(n135), .A2(n34), .ZN(n35) );
  NAND2_X1 U81 ( .A1(n123), .A2(n20), .ZN(n21) );
  AND2_X1 U82 ( .A1(n194), .A2(n104), .ZN(n102) );
  INV_X1 U83 ( .A(GE), .ZN(LT) );
  INV_X1 U84 ( .A(n93), .ZN(n186) );
  INV_X1 U85 ( .A(n79), .ZN(n174) );
  INV_X1 U86 ( .A(n65), .ZN(n162) );
  INV_X1 U87 ( .A(n51), .ZN(n150) );
  INV_X1 U88 ( .A(n37), .ZN(n138) );
  INV_X1 U89 ( .A(n23), .ZN(n126) );
  INV_X1 U90 ( .A(n90), .ZN(n89) );
  INV_X1 U91 ( .A(n76), .ZN(n75) );
  INV_X1 U92 ( .A(n62), .ZN(n61) );
  INV_X1 U93 ( .A(n48), .ZN(n47) );
  INV_X1 U94 ( .A(n34), .ZN(n33) );
  INV_X1 U95 ( .A(n20), .ZN(n19) );
  INV_X1 U96 ( .A(n104), .ZN(n103) );
  AOI21_X1 U97 ( .B1(n1), .B2(n2), .A(n3), .ZN(GE) );
  INV_X1 U98 ( .A(n4), .ZN(n2) );
  AOI22_X1 U99 ( .A1(B[30]), .A2(n5), .B1(n6), .B2(n7), .ZN(n4) );
  INV_X1 U100 ( .A(A[30]), .ZN(n5) );
  OAI21_X1 U101 ( .B1(n3), .B2(n109), .A(n1), .ZN(GT) );
  AOI22_X1 U102 ( .A1(A[30]), .A2(n111), .B1(n112), .B2(n7), .ZN(n109) );
  AOI21_X1 U103 ( .B1(n113), .B2(n114), .A(n115), .ZN(n112) );
  INV_X1 U104 ( .A(n9), .ZN(n115) );
  AOI22_X1 U105 ( .A1(n105), .A2(n106), .B1(A[1]), .B2(n107), .ZN(n101) );
  OR2_X1 U106 ( .A1(n107), .A2(A[1]), .ZN(n105) );
  NAND2_X1 U107 ( .A1(B[0]), .A2(n108), .ZN(n107) );
  NOR2_X1 U108 ( .A1(n108), .A2(B[0]), .ZN(n196) );
  NOR2_X1 U109 ( .A1(n191), .A2(B[4]), .ZN(n190) );
  NOR2_X1 U110 ( .A1(n180), .A2(B[8]), .ZN(n179) );
  NOR2_X1 U111 ( .A1(n168), .A2(B[12]), .ZN(n167) );
  NOR2_X1 U112 ( .A1(n156), .A2(B[16]), .ZN(n155) );
  NOR2_X1 U113 ( .A1(n144), .A2(B[20]), .ZN(n143) );
  NOR2_X1 U114 ( .A1(n132), .A2(B[24]), .ZN(n131) );
  NOR2_X1 U115 ( .A1(n120), .A2(B[28]), .ZN(n119) );
  NOR2_X1 U116 ( .A1(n187), .A2(B[5]), .ZN(n94) );
  NOR2_X1 U117 ( .A1(n175), .A2(B[9]), .ZN(n80) );
  NOR2_X1 U118 ( .A1(n163), .A2(B[13]), .ZN(n66) );
  NOR2_X1 U119 ( .A1(n151), .A2(B[17]), .ZN(n52) );
  NOR2_X1 U120 ( .A1(n139), .A2(B[21]), .ZN(n38) );
  NOR2_X1 U121 ( .A1(n127), .A2(B[25]), .ZN(n24) );
  NOR2_X1 U122 ( .A1(n116), .A2(B[29]), .ZN(n10) );
  NOR2_X1 U123 ( .A1(n192), .A2(B[3]), .ZN(n100) );
  NOR2_X1 U124 ( .A1(n181), .A2(B[7]), .ZN(n86) );
  NOR2_X1 U125 ( .A1(n169), .A2(B[11]), .ZN(n72) );
  NOR2_X1 U126 ( .A1(n157), .A2(B[15]), .ZN(n58) );
  NOR2_X1 U127 ( .A1(n145), .A2(B[19]), .ZN(n44) );
  NOR2_X1 U128 ( .A1(n133), .A2(B[23]), .ZN(n30) );
  NOR2_X1 U129 ( .A1(n121), .A2(B[27]), .ZN(n16) );
  NOR2_X1 U130 ( .A1(n110), .A2(A[31]), .ZN(n3) );
  INV_X1 U131 ( .A(n100), .ZN(n193) );
  OAI211_X1 U132 ( .C1(A[1]), .C2(n196), .A(n197), .B(n102), .ZN(n195) );
  NAND2_X1 U133 ( .A1(B[7]), .A2(n181), .ZN(n85) );
  NAND2_X1 U134 ( .A1(B[11]), .A2(n169), .ZN(n71) );
  NAND2_X1 U135 ( .A1(B[15]), .A2(n157), .ZN(n57) );
  NAND2_X1 U136 ( .A1(B[19]), .A2(n145), .ZN(n43) );
  NAND2_X1 U137 ( .A1(B[23]), .A2(n133), .ZN(n29) );
  NAND2_X1 U138 ( .A1(B[27]), .A2(n121), .ZN(n15) );
  NAND2_X1 U139 ( .A1(B[5]), .A2(n187), .ZN(n93) );
  NAND2_X1 U140 ( .A1(B[9]), .A2(n175), .ZN(n79) );
  NAND2_X1 U141 ( .A1(B[13]), .A2(n163), .ZN(n65) );
  NAND2_X1 U142 ( .A1(B[17]), .A2(n151), .ZN(n51) );
  NAND2_X1 U143 ( .A1(B[21]), .A2(n139), .ZN(n37) );
  NAND2_X1 U144 ( .A1(B[25]), .A2(n127), .ZN(n23) );
  NAND2_X1 U145 ( .A1(B[29]), .A2(n116), .ZN(n9) );
  NAND2_X1 U146 ( .A1(B[6]), .A2(n188), .ZN(n90) );
  NAND2_X1 U147 ( .A1(B[10]), .A2(n176), .ZN(n76) );
  NAND2_X1 U148 ( .A1(B[14]), .A2(n164), .ZN(n62) );
  NAND2_X1 U150 ( .A1(B[18]), .A2(n152), .ZN(n48) );
  NAND2_X1 U151 ( .A1(B[22]), .A2(n140), .ZN(n34) );
  NAND2_X1 U152 ( .A1(B[26]), .A2(n128), .ZN(n20) );
  NAND2_X1 U154 ( .A1(A[31]), .A2(n110), .ZN(n1) );
  AND2_X1 U155 ( .A1(B[4]), .A2(n191), .ZN(n97) );
  AND2_X1 U156 ( .A1(B[8]), .A2(n180), .ZN(n83) );
  AND2_X1 U157 ( .A1(B[12]), .A2(n168), .ZN(n69) );
  AND2_X1 U158 ( .A1(B[16]), .A2(n156), .ZN(n55) );
  AND2_X1 U159 ( .A1(B[20]), .A2(n144), .ZN(n41) );
  AND2_X1 U160 ( .A1(B[24]), .A2(n132), .ZN(n27) );
  AND2_X1 U161 ( .A1(B[28]), .A2(n120), .ZN(n13) );
  NAND2_X1 U162 ( .A1(B[3]), .A2(n192), .ZN(n99) );
  NAND2_X1 U163 ( .A1(B[2]), .A2(n198), .ZN(n104) );
  OR2_X1 U164 ( .A1(n188), .A2(B[6]), .ZN(n183) );
  OR2_X1 U165 ( .A1(n176), .A2(B[10]), .ZN(n171) );
  OR2_X1 U166 ( .A1(n164), .A2(B[14]), .ZN(n159) );
  OR2_X1 U167 ( .A1(n152), .A2(B[18]), .ZN(n147) );
  OR2_X1 U168 ( .A1(n140), .A2(B[22]), .ZN(n135) );
  OR2_X1 U169 ( .A1(n128), .A2(B[26]), .ZN(n123) );
  INV_X1 U170 ( .A(A[0]), .ZN(n108) );
  INV_X1 U171 ( .A(A[3]), .ZN(n192) );
  INV_X1 U172 ( .A(A[5]), .ZN(n187) );
  INV_X1 U173 ( .A(A[7]), .ZN(n181) );
  INV_X1 U174 ( .A(A[9]), .ZN(n175) );
  INV_X1 U175 ( .A(A[11]), .ZN(n169) );
  INV_X1 U176 ( .A(A[13]), .ZN(n163) );
  INV_X1 U177 ( .A(A[15]), .ZN(n157) );
  INV_X1 U178 ( .A(A[17]), .ZN(n151) );
  INV_X1 U179 ( .A(A[19]), .ZN(n145) );
  INV_X1 U180 ( .A(A[21]), .ZN(n139) );
  INV_X1 U181 ( .A(A[23]), .ZN(n133) );
  INV_X1 U182 ( .A(A[25]), .ZN(n127) );
  INV_X1 U183 ( .A(A[27]), .ZN(n121) );
  INV_X1 U184 ( .A(A[29]), .ZN(n116) );
  INV_X1 U185 ( .A(B[31]), .ZN(n110) );
  INV_X1 U186 ( .A(B[1]), .ZN(n106) );
  INV_X1 U187 ( .A(B[30]), .ZN(n111) );
  INV_X1 U188 ( .A(A[2]), .ZN(n198) );
  INV_X1 U189 ( .A(A[6]), .ZN(n188) );
  INV_X1 U190 ( .A(A[10]), .ZN(n176) );
  INV_X1 U191 ( .A(A[14]), .ZN(n164) );
  INV_X1 U192 ( .A(A[18]), .ZN(n152) );
  INV_X1 U193 ( .A(A[22]), .ZN(n140) );
  INV_X1 U194 ( .A(A[26]), .ZN(n128) );
  OR2_X1 U195 ( .A1(n198), .A2(B[2]), .ZN(n194) );
  INV_X1 U196 ( .A(A[4]), .ZN(n191) );
  INV_X1 U197 ( .A(A[8]), .ZN(n180) );
  INV_X1 U198 ( .A(A[12]), .ZN(n168) );
  INV_X1 U199 ( .A(A[16]), .ZN(n156) );
  INV_X1 U200 ( .A(A[20]), .ZN(n144) );
  INV_X1 U201 ( .A(A[24]), .ZN(n132) );
  INV_X1 U202 ( .A(A[28]), .ZN(n120) );
  INV_X1 U203 ( .A(n199), .ZN(n197) );
  AOI21_X1 U204 ( .B1(A[1]), .B2(n196), .A(n106), .ZN(n199) );
endmodule


module ALU_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200;

  NAND3_X1 U25 ( .A1(n72), .A2(n73), .A3(n74), .ZN(n69) );
  NAND3_X1 U26 ( .A1(n75), .A2(n76), .A3(n77), .ZN(n72) );
  XOR2_X1 U43 ( .A(n100), .B(B[30]), .Z(n8) );
  INV_X1 U1 ( .A(n60), .ZN(n168) );
  INV_X1 U2 ( .A(n40), .ZN(n140) );
  INV_X1 U3 ( .A(n20), .ZN(n112) );
  INV_X1 U4 ( .A(LT), .ZN(GE) );
  AOI211_X1 U5 ( .C1(n68), .C2(n69), .A(n70), .B(n71), .ZN(n62) );
  NOR2_X1 U6 ( .A1(n84), .A2(n85), .ZN(n68) );
  AOI211_X1 U7 ( .C1(n58), .C2(n59), .A(n60), .B(n61), .ZN(n52) );
  NOR2_X1 U8 ( .A1(n86), .A2(n87), .ZN(n58) );
  OAI211_X1 U9 ( .C1(n62), .C2(n63), .A(n64), .B(n65), .ZN(n59) );
  NAND2_X1 U10 ( .A1(n66), .A2(n67), .ZN(n63) );
  AOI211_X1 U11 ( .C1(n48), .C2(n49), .A(n50), .B(n51), .ZN(n42) );
  NOR2_X1 U12 ( .A1(n88), .A2(n89), .ZN(n48) );
  OAI211_X1 U13 ( .C1(n52), .C2(n53), .A(n54), .B(n55), .ZN(n49) );
  NAND2_X1 U14 ( .A1(n56), .A2(n57), .ZN(n53) );
  AOI211_X1 U15 ( .C1(n38), .C2(n39), .A(n40), .B(n41), .ZN(n32) );
  NOR2_X1 U16 ( .A1(n90), .A2(n91), .ZN(n38) );
  OAI211_X1 U17 ( .C1(n42), .C2(n43), .A(n44), .B(n45), .ZN(n39) );
  NAND2_X1 U18 ( .A1(n46), .A2(n47), .ZN(n43) );
  AOI211_X1 U19 ( .C1(n28), .C2(n29), .A(n30), .B(n31), .ZN(n22) );
  NOR2_X1 U20 ( .A1(n92), .A2(n93), .ZN(n28) );
  OAI211_X1 U21 ( .C1(n32), .C2(n33), .A(n34), .B(n35), .ZN(n29) );
  NAND2_X1 U22 ( .A1(n36), .A2(n37), .ZN(n33) );
  AOI211_X1 U23 ( .C1(n18), .C2(n19), .A(n20), .B(n21), .ZN(n12) );
  NOR2_X1 U24 ( .A1(n94), .A2(n95), .ZN(n18) );
  OAI211_X1 U27 ( .C1(n22), .C2(n23), .A(n24), .B(n25), .ZN(n19) );
  NAND2_X1 U28 ( .A1(n26), .A2(n27), .ZN(n23) );
  NOR2_X1 U29 ( .A1(n195), .A2(n196), .ZN(n80) );
  INV_X1 U30 ( .A(n76), .ZN(n196) );
  NOR2_X1 U31 ( .A1(n176), .A2(n86), .ZN(n65) );
  NOR2_X1 U32 ( .A1(n162), .A2(n88), .ZN(n55) );
  NOR2_X1 U33 ( .A1(n148), .A2(n90), .ZN(n45) );
  NOR2_X1 U34 ( .A1(n134), .A2(n92), .ZN(n35) );
  NOR2_X1 U35 ( .A1(n120), .A2(n94), .ZN(n25) );
  NOR2_X1 U36 ( .A1(n106), .A2(n96), .ZN(n15) );
  AOI21_X1 U37 ( .B1(n172), .B2(n173), .A(n87), .ZN(n167) );
  INV_X1 U38 ( .A(n61), .ZN(n173) );
  AOI21_X1 U39 ( .B1(n175), .B2(n65), .A(n176), .ZN(n172) );
  AOI21_X1 U40 ( .B1(n178), .B2(n64), .A(n179), .ZN(n175) );
  AOI21_X1 U41 ( .B1(n189), .B2(n74), .A(n190), .ZN(n186) );
  AOI21_X1 U42 ( .B1(n191), .B2(n73), .A(n192), .ZN(n189) );
  INV_X1 U44 ( .A(n75), .ZN(n192) );
  AOI21_X1 U45 ( .B1(n194), .B2(n80), .A(n195), .ZN(n191) );
  AOI21_X1 U46 ( .B1(n181), .B2(n182), .A(n183), .ZN(n178) );
  INV_X1 U47 ( .A(n70), .ZN(n182) );
  AOI21_X1 U48 ( .B1(n186), .B2(n187), .A(n85), .ZN(n181) );
  INV_X1 U49 ( .A(n71), .ZN(n187) );
  AOI21_X1 U50 ( .B1(n161), .B2(n55), .A(n162), .ZN(n158) );
  AOI21_X1 U51 ( .B1(n164), .B2(n54), .A(n165), .ZN(n161) );
  INV_X1 U52 ( .A(n56), .ZN(n165) );
  AOI21_X1 U53 ( .B1(n167), .B2(n168), .A(n169), .ZN(n164) );
  AOI21_X1 U54 ( .B1(n116), .B2(n117), .A(n95), .ZN(n111) );
  INV_X1 U55 ( .A(n21), .ZN(n117) );
  AOI21_X1 U56 ( .B1(n119), .B2(n25), .A(n120), .ZN(n116) );
  AOI21_X1 U57 ( .B1(n122), .B2(n24), .A(n123), .ZN(n119) );
  AOI21_X1 U58 ( .B1(n153), .B2(n154), .A(n155), .ZN(n150) );
  INV_X1 U59 ( .A(n50), .ZN(n154) );
  AOI21_X1 U60 ( .B1(n158), .B2(n159), .A(n89), .ZN(n153) );
  INV_X1 U61 ( .A(n51), .ZN(n159) );
  AOI21_X1 U62 ( .B1(n144), .B2(n145), .A(n91), .ZN(n139) );
  INV_X1 U63 ( .A(n41), .ZN(n145) );
  AOI21_X1 U64 ( .B1(n147), .B2(n45), .A(n148), .ZN(n144) );
  AOI21_X1 U65 ( .B1(n150), .B2(n44), .A(n151), .ZN(n147) );
  AOI21_X1 U66 ( .B1(n133), .B2(n35), .A(n134), .ZN(n130) );
  AOI21_X1 U67 ( .B1(n136), .B2(n34), .A(n137), .ZN(n133) );
  INV_X1 U68 ( .A(n36), .ZN(n137) );
  AOI21_X1 U69 ( .B1(n139), .B2(n140), .A(n141), .ZN(n136) );
  AOI21_X1 U70 ( .B1(n125), .B2(n126), .A(n127), .ZN(n122) );
  INV_X1 U71 ( .A(n30), .ZN(n126) );
  AOI21_X1 U72 ( .B1(n130), .B2(n131), .A(n93), .ZN(n125) );
  INV_X1 U73 ( .A(n31), .ZN(n131) );
  AOI21_X1 U74 ( .B1(n105), .B2(n15), .A(n106), .ZN(n102) );
  AOI21_X1 U75 ( .B1(n108), .B2(n14), .A(n109), .ZN(n105) );
  INV_X1 U76 ( .A(n16), .ZN(n109) );
  AOI21_X1 U77 ( .B1(n111), .B2(n112), .A(n113), .ZN(n108) );
  AOI21_X1 U78 ( .B1(n9), .B2(n10), .A(n11), .ZN(n7) );
  NOR2_X1 U79 ( .A1(n96), .A2(n97), .ZN(n9) );
  OAI211_X1 U80 ( .C1(n12), .C2(n13), .A(n14), .B(n15), .ZN(n10) );
  NAND2_X1 U81 ( .A1(n16), .A2(n17), .ZN(n13) );
  NOR2_X1 U82 ( .A1(n190), .A2(n84), .ZN(n74) );
  NAND2_X1 U83 ( .A1(n184), .A2(n67), .ZN(n70) );
  INV_X1 U84 ( .A(n183), .ZN(n184) );
  NAND2_X1 U85 ( .A1(n170), .A2(n57), .ZN(n60) );
  INV_X1 U86 ( .A(n169), .ZN(n170) );
  NAND2_X1 U87 ( .A1(n156), .A2(n47), .ZN(n50) );
  INV_X1 U88 ( .A(n155), .ZN(n156) );
  NAND2_X1 U89 ( .A1(n142), .A2(n37), .ZN(n40) );
  INV_X1 U90 ( .A(n141), .ZN(n142) );
  NAND2_X1 U91 ( .A1(n128), .A2(n27), .ZN(n30) );
  INV_X1 U92 ( .A(n127), .ZN(n128) );
  NAND2_X1 U93 ( .A1(n114), .A2(n17), .ZN(n20) );
  INV_X1 U94 ( .A(n113), .ZN(n114) );
  INV_X1 U95 ( .A(LE), .ZN(GT) );
  INV_X1 U96 ( .A(n66), .ZN(n179) );
  INV_X1 U97 ( .A(n46), .ZN(n151) );
  INV_X1 U98 ( .A(n26), .ZN(n123) );
  AOI21_X1 U99 ( .B1(n2), .B2(n3), .A(n4), .ZN(LE) );
  INV_X1 U100 ( .A(n5), .ZN(n3) );
  AOI22_X1 U101 ( .A1(A[30]), .A2(n6), .B1(n7), .B2(n8), .ZN(n5) );
  INV_X1 U102 ( .A(B[30]), .ZN(n6) );
  OAI21_X1 U103 ( .B1(n4), .B2(n98), .A(n2), .ZN(LT) );
  AOI22_X1 U104 ( .A1(B[30]), .A2(n100), .B1(n101), .B2(n8), .ZN(n98) );
  AOI21_X1 U105 ( .B1(n102), .B2(n103), .A(n97), .ZN(n101) );
  INV_X1 U106 ( .A(n11), .ZN(n103) );
  NOR2_X1 U107 ( .A1(n188), .A2(A[5]), .ZN(n71) );
  NOR2_X1 U108 ( .A1(n174), .A2(A[9]), .ZN(n61) );
  NOR2_X1 U109 ( .A1(n160), .A2(A[13]), .ZN(n51) );
  NOR2_X1 U110 ( .A1(n146), .A2(A[17]), .ZN(n41) );
  NOR2_X1 U111 ( .A1(n132), .A2(A[21]), .ZN(n31) );
  NOR2_X1 U112 ( .A1(n118), .A2(A[25]), .ZN(n21) );
  NOR2_X1 U113 ( .A1(n197), .A2(A[2]), .ZN(n195) );
  NOR2_X1 U114 ( .A1(n1), .A2(A[4]), .ZN(n190) );
  NOR2_X1 U115 ( .A1(n177), .A2(A[8]), .ZN(n176) );
  NOR2_X1 U116 ( .A1(n163), .A2(A[12]), .ZN(n162) );
  NOR2_X1 U117 ( .A1(n149), .A2(A[16]), .ZN(n148) );
  NOR2_X1 U118 ( .A1(n135), .A2(A[20]), .ZN(n134) );
  NOR2_X1 U119 ( .A1(n121), .A2(A[24]), .ZN(n120) );
  NOR2_X1 U120 ( .A1(n107), .A2(A[28]), .ZN(n106) );
  NOR2_X1 U121 ( .A1(n185), .A2(A[6]), .ZN(n183) );
  NOR2_X1 U122 ( .A1(n171), .A2(A[10]), .ZN(n169) );
  NOR2_X1 U123 ( .A1(n157), .A2(A[14]), .ZN(n155) );
  NOR2_X1 U124 ( .A1(n143), .A2(A[18]), .ZN(n141) );
  NOR2_X1 U125 ( .A1(n129), .A2(A[22]), .ZN(n127) );
  NOR2_X1 U126 ( .A1(n115), .A2(A[26]), .ZN(n113) );
  NOR2_X1 U127 ( .A1(n104), .A2(A[29]), .ZN(n11) );
  NOR2_X1 U128 ( .A1(n99), .A2(A[31]), .ZN(n4) );
  OAI211_X1 U129 ( .C1(A[1]), .C2(n78), .A(n79), .B(n80), .ZN(n77) );
  INV_X1 U130 ( .A(n82), .ZN(n78) );
  OAI21_X1 U131 ( .B1(n81), .B2(n82), .A(B[1]), .ZN(n79) );
  NAND2_X1 U132 ( .A1(A[0]), .A2(n83), .ZN(n82) );
  NAND2_X1 U133 ( .A1(A[6]), .A2(n185), .ZN(n67) );
  NAND2_X1 U134 ( .A1(A[10]), .A2(n171), .ZN(n57) );
  NAND2_X1 U135 ( .A1(A[14]), .A2(n157), .ZN(n47) );
  NAND2_X1 U136 ( .A1(A[18]), .A2(n143), .ZN(n37) );
  NAND2_X1 U137 ( .A1(A[22]), .A2(n129), .ZN(n27) );
  NAND2_X1 U138 ( .A1(A[26]), .A2(n115), .ZN(n17) );
  NAND2_X1 U139 ( .A1(A[31]), .A2(n99), .ZN(n2) );
  NAND2_X1 U140 ( .A1(A[7]), .A2(n180), .ZN(n66) );
  NAND2_X1 U141 ( .A1(A[11]), .A2(n166), .ZN(n56) );
  NAND2_X1 U142 ( .A1(A[15]), .A2(n152), .ZN(n46) );
  NAND2_X1 U143 ( .A1(A[19]), .A2(n138), .ZN(n36) );
  NAND2_X1 U144 ( .A1(A[23]), .A2(n124), .ZN(n26) );
  NAND2_X1 U145 ( .A1(A[27]), .A2(n110), .ZN(n16) );
  INV_X1 U146 ( .A(A[1]), .ZN(n81) );
  AND2_X1 U147 ( .A1(A[4]), .A2(n1), .ZN(n84) );
  AND2_X1 U148 ( .A1(A[8]), .A2(n177), .ZN(n86) );
  AND2_X1 U149 ( .A1(A[12]), .A2(n163), .ZN(n88) );
  AND2_X1 U150 ( .A1(A[16]), .A2(n149), .ZN(n90) );
  AND2_X1 U151 ( .A1(A[20]), .A2(n135), .ZN(n92) );
  AND2_X1 U152 ( .A1(A[24]), .A2(n121), .ZN(n94) );
  AND2_X1 U153 ( .A1(A[28]), .A2(n107), .ZN(n96) );
  AND2_X1 U154 ( .A1(A[5]), .A2(n188), .ZN(n85) );
  AND2_X1 U155 ( .A1(A[9]), .A2(n174), .ZN(n87) );
  AND2_X1 U156 ( .A1(A[13]), .A2(n160), .ZN(n89) );
  AND2_X1 U157 ( .A1(A[17]), .A2(n146), .ZN(n91) );
  AND2_X1 U158 ( .A1(A[21]), .A2(n132), .ZN(n93) );
  AND2_X1 U159 ( .A1(A[25]), .A2(n118), .ZN(n95) );
  AND2_X1 U160 ( .A1(A[29]), .A2(n104), .ZN(n97) );
  OR2_X1 U161 ( .A1(n180), .A2(A[7]), .ZN(n64) );
  OR2_X1 U162 ( .A1(n166), .A2(A[11]), .ZN(n54) );
  OR2_X1 U163 ( .A1(n152), .A2(A[15]), .ZN(n44) );
  OR2_X1 U164 ( .A1(n138), .A2(A[19]), .ZN(n34) );
  OR2_X1 U165 ( .A1(n124), .A2(A[23]), .ZN(n24) );
  OR2_X1 U166 ( .A1(n110), .A2(A[27]), .ZN(n14) );
  NAND2_X1 U167 ( .A1(A[2]), .A2(n197), .ZN(n76) );
  NAND2_X1 U168 ( .A1(A[3]), .A2(n193), .ZN(n75) );
  INV_X1 U169 ( .A(B[2]), .ZN(n197) );
  INV_X1 U170 ( .A(B[6]), .ZN(n185) );
  INV_X1 U171 ( .A(B[10]), .ZN(n171) );
  INV_X1 U172 ( .A(B[14]), .ZN(n157) );
  INV_X1 U173 ( .A(B[0]), .ZN(n83) );
  INV_X1 U174 ( .A(B[18]), .ZN(n143) );
  INV_X1 U175 ( .A(B[22]), .ZN(n129) );
  INV_X1 U176 ( .A(B[26]), .ZN(n115) );
  INV_X1 U177 ( .A(B[31]), .ZN(n99) );
  OR2_X1 U178 ( .A1(n193), .A2(A[3]), .ZN(n73) );
  INV_X1 U179 ( .A(A[30]), .ZN(n100) );
  INV_X1 U180 ( .A(B[3]), .ZN(n193) );
  INV_X1 U181 ( .A(B[7]), .ZN(n180) );
  INV_X1 U182 ( .A(B[11]), .ZN(n166) );
  INV_X1 U183 ( .A(B[15]), .ZN(n152) );
  INV_X1 U184 ( .A(B[19]), .ZN(n138) );
  INV_X1 U185 ( .A(B[23]), .ZN(n124) );
  INV_X1 U186 ( .A(B[27]), .ZN(n110) );
  INV_X1 U187 ( .A(B[4]), .ZN(n1) );
  INV_X1 U188 ( .A(B[5]), .ZN(n188) );
  INV_X1 U189 ( .A(B[8]), .ZN(n177) );
  INV_X1 U190 ( .A(B[9]), .ZN(n174) );
  INV_X1 U191 ( .A(B[12]), .ZN(n163) );
  INV_X1 U192 ( .A(B[13]), .ZN(n160) );
  INV_X1 U193 ( .A(B[16]), .ZN(n149) );
  INV_X1 U194 ( .A(B[17]), .ZN(n146) );
  INV_X1 U195 ( .A(B[20]), .ZN(n135) );
  INV_X1 U196 ( .A(B[21]), .ZN(n132) );
  INV_X1 U197 ( .A(B[24]), .ZN(n121) );
  INV_X1 U198 ( .A(B[25]), .ZN(n118) );
  INV_X1 U199 ( .A(B[28]), .ZN(n107) );
  INV_X1 U200 ( .A(B[29]), .ZN(n104) );
  INV_X1 U201 ( .A(n198), .ZN(n194) );
  OAI22_X1 U202 ( .A1(n199), .A2(B[1]), .B1(n81), .B2(n200), .ZN(n198) );
  AND2_X1 U203 ( .A1(n200), .A2(n81), .ZN(n199) );
  NOR2_X1 U204 ( .A1(n83), .A2(A[0]), .ZN(n200) );
endmodule


module ALU_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] ;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(\carry[31] ), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
endmodule


module ALU_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] ;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(\carry[31] ), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
endmodule


module ALU_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] , \B_not[31] , \B_not[30] , \B_not[29] , \B_not[28] ,
         \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] , \B_not[23] ,
         \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] , \B_not[18] ,
         \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] , \B_not[13] ,
         \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] , \B_not[8] ,
         \B_not[7] , \B_not[6] , \B_not[5] , \B_not[3] , \B_not[2] ,
         \B_not[1] , \B_not[0] , n1;

  FA_X1 U2_31 ( .A(A[31]), .B(\B_not[31] ), .CI(\carry[31] ), .S(DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(\B_not[30] ), .CI(\carry[30] ), .CO(\carry[31] ), 
        .S(DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(\B_not[29] ), .CI(\carry[29] ), .CO(\carry[30] ), 
        .S(DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(\B_not[28] ), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(\B_not[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(\B_not[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(\B_not[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(\B_not[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(\B_not[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(\B_not[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(\B_not[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(\B_not[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(\B_not[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(\B_not[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(\B_not[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(\B_not[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(\B_not[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(\B_not[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(\B_not[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(\B_not[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(\B_not[9] ), .CI(\carry[9] ), .CO(\carry[10] ), 
        .S(DIFF[9]) );
  FA_X1 U2_8 ( .A(A[8]), .B(\B_not[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(\B_not[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(\B_not[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(\B_not[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n1), .CI(\carry[4] ), .CO(\carry[5] ), .S(DIFF[4])
         );
  FA_X1 U2_3 ( .A(A[3]), .B(\B_not[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(\B_not[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(\B_not[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        DIFF[1]) );
  XNOR2_X1 U1 ( .A(A[0]), .B(\B_not[0] ), .ZN(DIFF[0]) );
  INV_X1 U2 ( .A(B[1]), .ZN(\B_not[1] ) );
  OR2_X1 U3 ( .A1(\B_not[0] ), .A2(A[0]), .ZN(\carry[1] ) );
  INV_X1 U4 ( .A(B[2]), .ZN(\B_not[2] ) );
  INV_X1 U5 ( .A(B[3]), .ZN(\B_not[3] ) );
  INV_X1 U6 ( .A(B[4]), .ZN(n1) );
  INV_X1 U7 ( .A(B[5]), .ZN(\B_not[5] ) );
  INV_X1 U8 ( .A(B[6]), .ZN(\B_not[6] ) );
  INV_X1 U9 ( .A(B[7]), .ZN(\B_not[7] ) );
  INV_X1 U10 ( .A(B[8]), .ZN(\B_not[8] ) );
  INV_X1 U11 ( .A(B[9]), .ZN(\B_not[9] ) );
  INV_X1 U12 ( .A(B[10]), .ZN(\B_not[10] ) );
  INV_X1 U13 ( .A(B[11]), .ZN(\B_not[11] ) );
  INV_X1 U14 ( .A(B[12]), .ZN(\B_not[12] ) );
  INV_X1 U15 ( .A(B[13]), .ZN(\B_not[13] ) );
  INV_X1 U16 ( .A(B[14]), .ZN(\B_not[14] ) );
  INV_X1 U17 ( .A(B[15]), .ZN(\B_not[15] ) );
  INV_X1 U18 ( .A(B[16]), .ZN(\B_not[16] ) );
  INV_X1 U19 ( .A(B[17]), .ZN(\B_not[17] ) );
  INV_X1 U20 ( .A(B[18]), .ZN(\B_not[18] ) );
  INV_X1 U21 ( .A(B[19]), .ZN(\B_not[19] ) );
  INV_X1 U22 ( .A(B[20]), .ZN(\B_not[20] ) );
  INV_X1 U23 ( .A(B[21]), .ZN(\B_not[21] ) );
  INV_X1 U24 ( .A(B[22]), .ZN(\B_not[22] ) );
  INV_X1 U25 ( .A(B[23]), .ZN(\B_not[23] ) );
  INV_X1 U26 ( .A(B[24]), .ZN(\B_not[24] ) );
  INV_X1 U27 ( .A(B[25]), .ZN(\B_not[25] ) );
  INV_X1 U28 ( .A(B[26]), .ZN(\B_not[26] ) );
  INV_X1 U29 ( .A(B[27]), .ZN(\B_not[27] ) );
  INV_X1 U30 ( .A(B[28]), .ZN(\B_not[28] ) );
  INV_X1 U31 ( .A(B[29]), .ZN(\B_not[29] ) );
  INV_X1 U32 ( .A(B[30]), .ZN(\B_not[30] ) );
  INV_X1 U33 ( .A(B[0]), .ZN(\B_not[0] ) );
  INV_X1 U34 ( .A(B[31]), .ZN(\B_not[31] ) );
endmodule


module ALU_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] , \B_not[31] , \B_not[30] , \B_not[29] , \B_not[28] ,
         \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] , \B_not[23] ,
         \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] , \B_not[18] ,
         \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] , \B_not[13] ,
         \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] , \B_not[8] ,
         \B_not[7] , \B_not[6] , \B_not[5] , \B_not[3] , \B_not[2] ,
         \B_not[1] , \B_not[0] , n1;

  FA_X1 U2_31 ( .A(A[31]), .B(\B_not[31] ), .CI(\carry[31] ), .S(DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(\B_not[30] ), .CI(\carry[30] ), .CO(\carry[31] ), 
        .S(DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(\B_not[29] ), .CI(\carry[29] ), .CO(\carry[30] ), 
        .S(DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(\B_not[28] ), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(\B_not[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(\B_not[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(\B_not[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(\B_not[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(\B_not[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(\B_not[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(\B_not[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(\B_not[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(\B_not[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(\B_not[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(\B_not[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(\B_not[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(\B_not[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(\B_not[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(\B_not[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(\B_not[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(\B_not[9] ), .CI(\carry[9] ), .CO(\carry[10] ), 
        .S(DIFF[9]) );
  FA_X1 U2_8 ( .A(A[8]), .B(\B_not[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(\B_not[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(\B_not[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(\B_not[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n1), .CI(\carry[4] ), .CO(\carry[5] ), .S(DIFF[4])
         );
  FA_X1 U2_3 ( .A(A[3]), .B(\B_not[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(\B_not[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(\B_not[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        DIFF[1]) );
  XNOR2_X1 U1 ( .A(A[0]), .B(\B_not[0] ), .ZN(DIFF[0]) );
  INV_X1 U2 ( .A(B[13]), .ZN(\B_not[13] ) );
  INV_X1 U3 ( .A(B[14]), .ZN(\B_not[14] ) );
  INV_X1 U4 ( .A(B[1]), .ZN(\B_not[1] ) );
  OR2_X1 U5 ( .A1(\B_not[0] ), .A2(A[0]), .ZN(\carry[1] ) );
  INV_X1 U6 ( .A(B[2]), .ZN(\B_not[2] ) );
  INV_X1 U7 ( .A(B[3]), .ZN(\B_not[3] ) );
  INV_X1 U8 ( .A(B[4]), .ZN(n1) );
  INV_X1 U9 ( .A(B[5]), .ZN(\B_not[5] ) );
  INV_X1 U10 ( .A(B[6]), .ZN(\B_not[6] ) );
  INV_X1 U11 ( .A(B[7]), .ZN(\B_not[7] ) );
  INV_X1 U12 ( .A(B[8]), .ZN(\B_not[8] ) );
  INV_X1 U13 ( .A(B[9]), .ZN(\B_not[9] ) );
  INV_X1 U14 ( .A(B[10]), .ZN(\B_not[10] ) );
  INV_X1 U15 ( .A(B[11]), .ZN(\B_not[11] ) );
  INV_X1 U16 ( .A(B[12]), .ZN(\B_not[12] ) );
  INV_X1 U17 ( .A(B[15]), .ZN(\B_not[15] ) );
  INV_X1 U18 ( .A(B[16]), .ZN(\B_not[16] ) );
  INV_X1 U19 ( .A(B[17]), .ZN(\B_not[17] ) );
  INV_X1 U20 ( .A(B[18]), .ZN(\B_not[18] ) );
  INV_X1 U21 ( .A(B[19]), .ZN(\B_not[19] ) );
  INV_X1 U22 ( .A(B[20]), .ZN(\B_not[20] ) );
  INV_X1 U23 ( .A(B[21]), .ZN(\B_not[21] ) );
  INV_X1 U24 ( .A(B[22]), .ZN(\B_not[22] ) );
  INV_X1 U25 ( .A(B[23]), .ZN(\B_not[23] ) );
  INV_X1 U26 ( .A(B[24]), .ZN(\B_not[24] ) );
  INV_X1 U27 ( .A(B[25]), .ZN(\B_not[25] ) );
  INV_X1 U28 ( .A(B[26]), .ZN(\B_not[26] ) );
  INV_X1 U29 ( .A(B[27]), .ZN(\B_not[27] ) );
  INV_X1 U30 ( .A(B[28]), .ZN(\B_not[28] ) );
  INV_X1 U31 ( .A(B[29]), .ZN(\B_not[29] ) );
  INV_X1 U32 ( .A(B[30]), .ZN(\B_not[30] ) );
  INV_X1 U33 ( .A(B[0]), .ZN(\B_not[0] ) );
  INV_X1 U34 ( .A(B[31]), .ZN(\B_not[31] ) );
endmodule


module mmu_out_iram ( from_iram, flush, to_if_id_reg );
  input [31:0] from_iram;
  output [31:0] to_if_id_reg;
  input flush;
  wire   n2, n5, n6, n7;

  BUF_X1 U3 ( .A(n2), .Z(n6) );
  BUF_X1 U4 ( .A(n2), .Z(n5) );
  BUF_X1 U5 ( .A(n2), .Z(n7) );
  INV_X1 U6 ( .A(flush), .ZN(n2) );
  AND2_X1 U7 ( .A1(from_iram[0]), .A2(n7), .ZN(to_if_id_reg[0]) );
  AND2_X1 U8 ( .A1(from_iram[1]), .A2(n6), .ZN(to_if_id_reg[1]) );
  AND2_X1 U9 ( .A1(from_iram[2]), .A2(n5), .ZN(to_if_id_reg[2]) );
  AND2_X1 U10 ( .A1(from_iram[3]), .A2(n5), .ZN(to_if_id_reg[3]) );
  AND2_X1 U11 ( .A1(from_iram[4]), .A2(n5), .ZN(to_if_id_reg[4]) );
  AND2_X1 U12 ( .A1(from_iram[5]), .A2(n5), .ZN(to_if_id_reg[5]) );
  AND2_X1 U13 ( .A1(from_iram[6]), .A2(n5), .ZN(to_if_id_reg[6]) );
  AND2_X1 U14 ( .A1(from_iram[7]), .A2(n5), .ZN(to_if_id_reg[7]) );
  AND2_X1 U15 ( .A1(from_iram[8]), .A2(n5), .ZN(to_if_id_reg[8]) );
  AND2_X1 U16 ( .A1(from_iram[9]), .A2(n5), .ZN(to_if_id_reg[9]) );
  AND2_X1 U17 ( .A1(from_iram[10]), .A2(n7), .ZN(to_if_id_reg[10]) );
  AND2_X1 U18 ( .A1(from_iram[11]), .A2(n7), .ZN(to_if_id_reg[11]) );
  AND2_X1 U19 ( .A1(from_iram[12]), .A2(n7), .ZN(to_if_id_reg[12]) );
  AND2_X1 U20 ( .A1(from_iram[13]), .A2(n7), .ZN(to_if_id_reg[13]) );
  AND2_X1 U21 ( .A1(from_iram[14]), .A2(n6), .ZN(to_if_id_reg[14]) );
  AND2_X1 U22 ( .A1(from_iram[15]), .A2(n6), .ZN(to_if_id_reg[15]) );
  AND2_X1 U23 ( .A1(from_iram[16]), .A2(n6), .ZN(to_if_id_reg[16]) );
  AND2_X1 U24 ( .A1(from_iram[17]), .A2(n6), .ZN(to_if_id_reg[17]) );
  AND2_X1 U25 ( .A1(from_iram[18]), .A2(n6), .ZN(to_if_id_reg[18]) );
  AND2_X1 U26 ( .A1(from_iram[19]), .A2(n6), .ZN(to_if_id_reg[19]) );
  AND2_X1 U27 ( .A1(from_iram[20]), .A2(n6), .ZN(to_if_id_reg[20]) );
  AND2_X1 U28 ( .A1(from_iram[21]), .A2(n6), .ZN(to_if_id_reg[21]) );
  AND2_X1 U29 ( .A1(from_iram[22]), .A2(n6), .ZN(to_if_id_reg[22]) );
  AND2_X1 U30 ( .A1(from_iram[23]), .A2(n6), .ZN(to_if_id_reg[23]) );
  AND2_X1 U31 ( .A1(from_iram[24]), .A2(n6), .ZN(to_if_id_reg[24]) );
  AND2_X1 U32 ( .A1(from_iram[25]), .A2(n5), .ZN(to_if_id_reg[25]) );
  AND2_X1 U33 ( .A1(from_iram[27]), .A2(n5), .ZN(to_if_id_reg[27]) );
  AND2_X1 U34 ( .A1(from_iram[29]), .A2(n5), .ZN(to_if_id_reg[29]) );
  OR2_X1 U35 ( .A1(flush), .A2(from_iram[26]), .ZN(to_if_id_reg[26]) );
  OR2_X1 U36 ( .A1(flush), .A2(from_iram[28]), .ZN(to_if_id_reg[28]) );
  OR2_X1 U37 ( .A1(flush), .A2(from_iram[30]), .ZN(to_if_id_reg[30]) );
  AND2_X1 U38 ( .A1(from_iram[31]), .A2(n5), .ZN(to_if_id_reg[31]) );
endmodule


module mmu_in_iram ( from_pc, to_iram );
  input [31:0] from_pc;
  output [31:0] to_iram;
  wire   \from_pc[31] , \from_pc[30] , \from_pc[29] , \from_pc[28] ,
         \from_pc[27] , \from_pc[26] , \from_pc[25] , \from_pc[24] ,
         \from_pc[23] , \from_pc[22] , \from_pc[21] , \from_pc[20] ,
         \from_pc[19] , \from_pc[18] , \from_pc[17] , \from_pc[16] ,
         \from_pc[15] , \from_pc[14] , \from_pc[13] , \from_pc[12] ,
         \from_pc[11] , \from_pc[10] , \from_pc[9] , \from_pc[8] ,
         \from_pc[7] , \from_pc[6] , \from_pc[5] , \from_pc[4] , \from_pc[3] ,
         \from_pc[2] ;
  assign to_iram[31] = 1'b0;
  assign to_iram[30] = 1'b0;
  assign to_iram[29] = \from_pc[31] ;
  assign \from_pc[31]  = from_pc[31];
  assign to_iram[28] = \from_pc[30] ;
  assign \from_pc[30]  = from_pc[30];
  assign to_iram[27] = \from_pc[29] ;
  assign \from_pc[29]  = from_pc[29];
  assign to_iram[26] = \from_pc[28] ;
  assign \from_pc[28]  = from_pc[28];
  assign to_iram[25] = \from_pc[27] ;
  assign \from_pc[27]  = from_pc[27];
  assign to_iram[24] = \from_pc[26] ;
  assign \from_pc[26]  = from_pc[26];
  assign to_iram[23] = \from_pc[25] ;
  assign \from_pc[25]  = from_pc[25];
  assign to_iram[22] = \from_pc[24] ;
  assign \from_pc[24]  = from_pc[24];
  assign to_iram[21] = \from_pc[23] ;
  assign \from_pc[23]  = from_pc[23];
  assign to_iram[20] = \from_pc[22] ;
  assign \from_pc[22]  = from_pc[22];
  assign to_iram[19] = \from_pc[21] ;
  assign \from_pc[21]  = from_pc[21];
  assign to_iram[18] = \from_pc[20] ;
  assign \from_pc[20]  = from_pc[20];
  assign to_iram[17] = \from_pc[19] ;
  assign \from_pc[19]  = from_pc[19];
  assign to_iram[16] = \from_pc[18] ;
  assign \from_pc[18]  = from_pc[18];
  assign to_iram[15] = \from_pc[17] ;
  assign \from_pc[17]  = from_pc[17];
  assign to_iram[14] = \from_pc[16] ;
  assign \from_pc[16]  = from_pc[16];
  assign to_iram[13] = \from_pc[15] ;
  assign \from_pc[15]  = from_pc[15];
  assign to_iram[12] = \from_pc[14] ;
  assign \from_pc[14]  = from_pc[14];
  assign to_iram[11] = \from_pc[13] ;
  assign \from_pc[13]  = from_pc[13];
  assign to_iram[10] = \from_pc[12] ;
  assign \from_pc[12]  = from_pc[12];
  assign to_iram[9] = \from_pc[11] ;
  assign \from_pc[11]  = from_pc[11];
  assign to_iram[8] = \from_pc[10] ;
  assign \from_pc[10]  = from_pc[10];
  assign to_iram[7] = \from_pc[9] ;
  assign \from_pc[9]  = from_pc[9];
  assign to_iram[6] = \from_pc[8] ;
  assign \from_pc[8]  = from_pc[8];
  assign to_iram[5] = \from_pc[7] ;
  assign \from_pc[7]  = from_pc[7];
  assign to_iram[4] = \from_pc[6] ;
  assign \from_pc[6]  = from_pc[6];
  assign to_iram[3] = \from_pc[5] ;
  assign \from_pc[5]  = from_pc[5];
  assign to_iram[2] = \from_pc[4] ;
  assign \from_pc[4]  = from_pc[4];
  assign to_iram[1] = \from_pc[3] ;
  assign \from_pc[3]  = from_pc[3];
  assign to_iram[0] = \from_pc[2] ;
  assign \from_pc[2]  = from_pc[2];

endmodule


module increment_pc_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , n1;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X1 U3 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  XOR2_X1 U5 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  XOR2_X1 U7 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  XOR2_X1 U9 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  XOR2_X1 U11 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  XOR2_X1 U13 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  XOR2_X1 U15 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  XOR2_X1 U17 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  XOR2_X1 U19 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  XOR2_X1 U21 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X1 U25 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  XOR2_X1 U27 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  XOR2_X1 U29 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  XOR2_X1 U31 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  XOR2_X1 U33 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  XOR2_X1 U35 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  XOR2_X1 U37 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  XOR2_X1 U39 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  XOR2_X1 U41 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  XOR2_X1 U43 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  XOR2_X1 U45 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  XOR2_X1 U47 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  XOR2_X1 U49 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  XOR2_X1 U51 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  XOR2_X1 U53 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U55 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  XOR2_X1 U57 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  XNOR2_X1 U1 ( .A(A[31]), .B(n1), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n1) );
  AND2_X1 U4 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  AND2_X1 U6 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  AND2_X1 U8 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  AND2_X1 U10 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  AND2_X1 U12 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  AND2_X1 U14 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  AND2_X1 U16 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  AND2_X1 U18 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  AND2_X1 U20 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  AND2_X1 U22 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  AND2_X1 U24 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  AND2_X1 U26 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  AND2_X1 U28 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  AND2_X1 U30 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  AND2_X1 U32 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  AND2_X1 U34 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  AND2_X1 U36 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  AND2_X1 U38 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U40 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U42 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  AND2_X1 U44 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  AND2_X1 U46 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  AND2_X1 U48 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  AND2_X1 U50 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  AND2_X1 U52 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  AND2_X1 U54 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  AND2_X1 U56 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  INV_X1 U58 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module dram_block ( address, data_write, mem_op, Data_out, unaligned, 
        data_read, read_op, write_op, nibble, write_byte, Address_toRAM, 
        Data_in );
  input [31:0] address;
  input [31:0] data_write;
  input [5:0] mem_op;
  input [31:0] Data_out;
  output [31:0] data_read;
  output [1:0] nibble;
  output [31:0] Address_toRAM;
  output [31:0] Data_in;
  output unaligned, read_op, write_op, write_byte;

  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign Address_toRAM[31] = 1'b0;
  assign Address_toRAM[30] = 1'b0;

  mmu_in_dram mmu_in0 ( .mem_op(mem_op), .aligned_address(address), .data(
        data_write), .unaligned(unaligned), .nibble(nibble), .write_op(
        write_op), .read_op(read_op), .mem_address({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, Address_toRAM[29:0]}), .mem_data(Data_in), 
        .write_byte(write_byte) );
  mmu_out_dram mmu_out0 ( .data_ram(Data_out), .mem_op(mem_op), .nibble(nibble), .unaligned(unaligned), .data_read(data_read) );
endmodule


module ALU ( alu_op, a, b, ovf, zero, res );
  input [4:0] alu_op;
  input [31:0] a;
  input [31:0] b;
  output [31:0] res;
  output ovf, zero;
  wire   N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539,
         N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550,
         N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N629, N630, N631,
         N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N658, N659, N660, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, n694, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n715, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899;
  assign n694 = b[4];

  DLH_X1 ovf_reg ( .G(N766), .D(N767), .Q(ovf) );
  NOR2_X2 U567 ( .A1(n306), .A2(n357), .ZN(n191) );
  NAND3_X1 U713 ( .A1(n332), .A2(n333), .A3(n334), .ZN(res[31]) );
  NAND3_X1 U714 ( .A1(a[31]), .A2(n359), .A3(n472), .ZN(n471) );
  NAND3_X1 U715 ( .A1(n299), .A2(n736), .A3(n843), .ZN(n734) );
  OAI33_X1 U716 ( .A1(n790), .A2(alu_op[4]), .A3(n791), .B1(n792), .B2(n793), 
        .B3(n794), .ZN(n789) );
  OAI33_X1 U717 ( .A1(n833), .A2(b[31]), .A3(a[31]), .B1(n831), .B2(N560), 
        .B3(n712), .ZN(n832) );
  ALU_DW01_sub_0 sub_76 ( .A(a), .B({b[31:5], n694, b[3:0]}), .CI(1'b0), 
        .DIFF({N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, 
        N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, 
        N638, N637, N636, N635, N634, N633, N632, N631, N630, N629}) );
  ALU_DW01_sub_1 sub_67 ( .A(a), .B({b[31:5], n694, b[3:0]}), .CI(1'b0), 
        .DIFF({N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, 
        N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, 
        N603, N602, N601, N600, N599, N598, N597, N596, N595, N594}) );
  ALU_DW01_add_0 add_64 ( .A(a), .B({b[31:5], n694, b[3:0]}), .CI(1'b0), .SUM(
        {N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, 
        N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, 
        N570, N569, N568, N567, N566, N565, N564, N563, N562}) );
  ALU_DW01_add_1 add_60 ( .A(a), .B({b[31:5], n694, b[3:0]}), .CI(1'b0), .SUM(
        {N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, 
        N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, 
        N537, N536, N535, N534, N533, N532, N531, N530, N529}) );
  ALU_DW01_cmp6_0 r95 ( .A(a), .B({b[31:5], n694, b[3:0]}), .TC(1'b1), .LT(
        N759), .GT(N760), .LE(N761), .GE(N762) );
  ALU_DW01_cmp6_1 r94 ( .A(a), .B({b[31:5], n694, b[3:0]}), .TC(1'b0), .LT(
        N763), .GT(N764), .EQ(N757), .GE(N765), .NE(N758) );
  AOI221_X1 U6 ( .B1(n344), .B2(a[26]), .C1(n865), .C2(a[25]), .A(n815), .ZN(
        n521) );
  OAI222_X1 U7 ( .A1(n862), .A2(n609), .B1(n860), .B2(n774), .C1(n834), .C2(
        n401), .ZN(n274) );
  OAI221_X1 U8 ( .B1(n860), .B2(n304), .C1(n863), .C2(n290), .A(n779), .ZN(
        n275) );
  NOR2_X1 U9 ( .A1(n624), .A2(n737), .ZN(n310) );
  NOR2_X1 U10 ( .A1(n362), .A2(n694), .ZN(n472) );
  INV_X1 U11 ( .A(n321), .ZN(n200) );
  INV_X1 U14 ( .A(n735), .ZN(n695) );
  INV_X1 U15 ( .A(n898), .ZN(n894) );
  INV_X1 U16 ( .A(n897), .ZN(n895) );
  INV_X1 U17 ( .A(n887), .ZN(n886) );
  INV_X1 U18 ( .A(n889), .ZN(n888) );
  INV_X1 U19 ( .A(n898), .ZN(n896) );
  INV_X1 U20 ( .A(n198), .ZN(n230) );
  INV_X1 U21 ( .A(n899), .ZN(n893) );
  INV_X1 U22 ( .A(n892), .ZN(n890) );
  INV_X1 U23 ( .A(n892), .ZN(n891) );
  INV_X1 U24 ( .A(n191), .ZN(n229) );
  NAND2_X1 U25 ( .A1(n837), .A2(n592), .ZN(n321) );
  INV_X1 U26 ( .A(n208), .ZN(n225) );
  NOR2_X1 U27 ( .A1(n183), .A2(n359), .ZN(n682) );
  INV_X1 U28 ( .A(n487), .ZN(n468) );
  INV_X1 U29 ( .A(n715), .ZN(n885) );
  NOR2_X1 U30 ( .A1(n470), .A2(n839), .ZN(n735) );
  INV_X1 U31 ( .A(n206), .ZN(n232) );
  NAND2_X1 U32 ( .A1(n183), .A2(n752), .ZN(n299) );
  BUF_X1 U33 ( .A(n209), .Z(n880) );
  BUF_X1 U34 ( .A(n209), .Z(n879) );
  BUF_X1 U35 ( .A(n211), .Z(n873) );
  BUF_X1 U36 ( .A(n211), .Z(n874) );
  BUF_X1 U37 ( .A(n211), .Z(n875) );
  BUF_X1 U38 ( .A(n209), .Z(n881) );
  INV_X1 U39 ( .A(n372), .ZN(n361) );
  INV_X1 U40 ( .A(n841), .ZN(n359) );
  INV_X1 U41 ( .A(n852), .ZN(n357) );
  BUF_X1 U42 ( .A(n855), .Z(n859) );
  BUF_X1 U43 ( .A(n855), .Z(n858) );
  BUF_X1 U44 ( .A(n855), .Z(n857) );
  BUF_X1 U45 ( .A(n856), .Z(n860) );
  BUF_X1 U46 ( .A(n856), .Z(n861) );
  NOR2_X1 U47 ( .A1(n639), .A2(n306), .ZN(n487) );
  NOR2_X1 U48 ( .A1(n306), .A2(n461), .ZN(n198) );
  NAND2_X1 U49 ( .A1(n854), .A2(n592), .ZN(n206) );
  INV_X1 U50 ( .A(n279), .ZN(n193) );
  NOR4_X1 U51 ( .A1(res[16]), .A2(res[15]), .A3(res[14]), .A4(res[13]), .ZN(
        n167) );
  NOR2_X1 U52 ( .A1(n463), .A2(n359), .ZN(n369) );
  INV_X1 U53 ( .A(n309), .ZN(n470) );
  NAND2_X1 U54 ( .A1(n310), .A2(n592), .ZN(n208) );
  NAND2_X1 U55 ( .A1(n463), .A2(n458), .ZN(n592) );
  OAI22_X1 U56 ( .A1(n388), .A2(n715), .B1(n387), .B2(n229), .ZN(n697) );
  OAI22_X1 U57 ( .A1(n358), .A2(n715), .B1(n356), .B2(n229), .ZN(n676) );
  OAI22_X1 U58 ( .A1(n228), .A2(n229), .B1(n230), .B2(n231), .ZN(n227) );
  OAI22_X1 U59 ( .A1(n490), .A2(n752), .B1(n278), .B2(n206), .ZN(n780) );
  OAI22_X1 U60 ( .A1(n278), .A2(n321), .B1(n701), .B2(n206), .ZN(n700) );
  OAI22_X1 U61 ( .A1(n571), .A2(n468), .B1(n423), .B2(n230), .ZN(n656) );
  OAI22_X1 U62 ( .A1(n462), .A2(n468), .B1(n356), .B2(n230), .ZN(n630) );
  OAI22_X1 U63 ( .A1(n519), .A2(n468), .B1(n597), .B2(n230), .ZN(n596) );
  OAI22_X1 U64 ( .A1(n490), .A2(n463), .B1(n491), .B2(n230), .ZN(n489) );
  OAI22_X1 U65 ( .A1(n358), .A2(n468), .B1(n469), .B2(n230), .ZN(n467) );
  OAI22_X1 U66 ( .A1(n277), .A2(n206), .B1(n278), .B2(n279), .ZN(n276) );
  OAI22_X1 U67 ( .A1(n277), .A2(n321), .B1(n701), .B2(n279), .ZN(n775) );
  OAI22_X1 U68 ( .A1(n744), .A2(n321), .B1(n593), .B2(n279), .ZN(n743) );
  OAI22_X1 U69 ( .A1(n460), .A2(n468), .B1(n462), .B2(n230), .ZN(n675) );
  OAI22_X1 U70 ( .A1(n205), .A2(n279), .B1(n293), .B2(n208), .ZN(n292) );
  OAI22_X1 U71 ( .A1(n259), .A2(n206), .B1(n260), .B2(n208), .ZN(n258) );
  OAI22_X1 U72 ( .A1(n356), .A2(n715), .B1(n259), .B2(n321), .ZN(n761) );
  INV_X1 U73 ( .A(n221), .ZN(n183) );
  OR2_X1 U74 ( .A1(n306), .A2(n359), .ZN(n715) );
  INV_X1 U75 ( .A(n179), .ZN(n752) );
  AOI21_X1 U76 ( .B1(n432), .B2(n361), .A(n433), .ZN(n431) );
  INV_X1 U77 ( .A(n369), .ZN(n432) );
  INV_X1 U78 ( .A(n549), .ZN(n532) );
  INV_X1 U79 ( .A(n548), .ZN(n533) );
  NOR2_X1 U80 ( .A1(n343), .A2(n434), .ZN(n372) );
  OAI22_X1 U81 ( .A1(n462), .A2(n532), .B1(n460), .B2(n533), .ZN(n531) );
  BUF_X1 U82 ( .A(n203), .Z(n882) );
  BUF_X1 U83 ( .A(n203), .Z(n883) );
  BUF_X1 U84 ( .A(n210), .Z(n876) );
  BUF_X1 U85 ( .A(n210), .Z(n877) );
  NAND2_X1 U86 ( .A1(n179), .A2(n841), .ZN(n693) );
  BUF_X1 U87 ( .A(n210), .Z(n878) );
  BUF_X1 U88 ( .A(n203), .Z(n884) );
  INV_X1 U89 ( .A(n190), .ZN(n887) );
  INV_X1 U90 ( .A(n827), .ZN(n211) );
  INV_X1 U91 ( .A(n826), .ZN(n209) );
  INV_X1 U92 ( .A(n865), .ZN(n862) );
  INV_X1 U93 ( .A(n872), .ZN(n871) );
  INV_X1 U94 ( .A(n872), .ZN(n870) );
  INV_X1 U95 ( .A(n872), .ZN(n869) );
  INV_X1 U96 ( .A(n865), .ZN(n864) );
  INV_X1 U97 ( .A(n865), .ZN(n863) );
  OAI22_X1 U98 ( .A1(n540), .A2(n357), .B1(n541), .B2(n359), .ZN(n537) );
  INV_X1 U99 ( .A(n310), .ZN(n639) );
  OAI22_X1 U100 ( .A1(n423), .A2(n357), .B1(n424), .B2(n359), .ZN(n422) );
  OAI22_X1 U101 ( .A1(n387), .A2(n357), .B1(n388), .B2(n359), .ZN(n386) );
  OAI22_X1 U102 ( .A1(n356), .A2(n357), .B1(n358), .B2(n359), .ZN(n355) );
  OAI21_X1 U103 ( .B1(n576), .B2(n639), .A(n653), .ZN(n611) );
  OAI21_X1 U104 ( .B1(n580), .B2(n639), .A(n653), .ZN(n610) );
  OAI21_X1 U105 ( .B1(n576), .B2(n461), .A(n577), .ZN(n284) );
  INV_X1 U106 ( .A(n410), .ZN(n580) );
  INV_X1 U107 ( .A(n661), .ZN(n231) );
  INV_X1 U108 ( .A(n412), .ZN(n576) );
  BUF_X1 U109 ( .A(n326), .Z(n855) );
  OR2_X1 U110 ( .A1(n220), .A2(n503), .ZN(n217) );
  OR2_X1 U111 ( .A1(n537), .A2(n503), .ZN(n255) );
  NAND2_X1 U112 ( .A1(n826), .A2(n827), .ZN(N766) );
  BUF_X1 U113 ( .A(n326), .Z(n856) );
  NOR2_X1 U114 ( .A1(n362), .A2(n308), .ZN(n179) );
  NOR2_X1 U115 ( .A1(n308), .A2(n434), .ZN(n221) );
  NOR2_X1 U116 ( .A1(n752), .A2(n712), .ZN(n309) );
  NOR2_X1 U117 ( .A1(n478), .A2(n359), .ZN(n549) );
  AOI222_X1 U118 ( .A1(n191), .A2(n197), .B1(n200), .B2(n291), .C1(n232), .C2(
        n199), .ZN(n282) );
  AOI222_X1 U119 ( .A1(n193), .A2(n233), .B1(n309), .B2(n310), .C1(n225), .C2(
        n237), .ZN(n297) );
  AOI222_X1 U120 ( .A1(N563), .A2(n884), .B1(n225), .B2(n294), .C1(n885), .C2(
        n197), .ZN(n599) );
  NOR4_X1 U121 ( .A1(res[9]), .A2(res[8]), .A3(res[7]), .A4(res[6]), .ZN(n173)
         );
  NOR4_X1 U122 ( .A1(res[23]), .A2(res[22]), .A3(res[21]), .A4(res[20]), .ZN(
        n169) );
  NOR4_X1 U123 ( .A1(res[1]), .A2(res[19]), .A3(res[18]), .A4(res[17]), .ZN(
        n168) );
  AOI221_X1 U124 ( .B1(n452), .B2(n514), .C1(n515), .C2(n220), .A(n516), .ZN(
        n513) );
  OAI222_X1 U125 ( .A1(n519), .A2(n359), .B1(n228), .B2(n357), .C1(n461), .C2(
        n231), .ZN(n514) );
  OAI21_X1 U126 ( .B1(n517), .B2(n485), .A(n470), .ZN(n516) );
  INV_X1 U127 ( .A(n518), .ZN(n517) );
  AOI221_X1 U128 ( .B1(n191), .B2(n192), .C1(n193), .C2(n194), .A(n195), .ZN(
        n176) );
  INV_X1 U129 ( .A(n196), .ZN(n195) );
  AOI22_X1 U130 ( .A1(n197), .A2(n198), .B1(n199), .B2(n200), .ZN(n196) );
  AOI221_X1 U131 ( .B1(n193), .B2(n626), .C1(n200), .C2(n254), .A(n685), .ZN(
        n672) );
  OAI22_X1 U132 ( .A1(n540), .A2(n208), .B1(n260), .B2(n206), .ZN(n685) );
  AOI221_X1 U133 ( .B1(n487), .B2(n483), .C1(N584), .C2(n883), .A(n564), .ZN(
        n545) );
  OAI22_X1 U134 ( .A1(n388), .A2(n230), .B1(n491), .B2(n229), .ZN(n564) );
  AOI221_X1 U135 ( .B1(n487), .B2(n202), .C1(N583), .C2(n883), .A(n582), .ZN(
        n566) );
  OAI22_X1 U136 ( .A1(n424), .A2(n230), .B1(n508), .B2(n229), .ZN(n582) );
  AOI221_X1 U137 ( .B1(n232), .B2(n233), .C1(N570), .C2(n882), .A(n234), .ZN(
        n213) );
  INV_X1 U138 ( .A(n235), .ZN(n234) );
  AOI22_X1 U139 ( .A1(n236), .A2(n200), .B1(n237), .B2(n193), .ZN(n235) );
  AOI221_X1 U140 ( .B1(n487), .B2(n542), .C1(N585), .C2(n883), .A(n543), .ZN(
        n527) );
  OAI22_X1 U141 ( .A1(n358), .A2(n230), .B1(n469), .B2(n229), .ZN(n543) );
  NOR4_X1 U142 ( .A1(res[12]), .A2(res[11]), .A3(res[10]), .A4(res[0]), .ZN(
        n166) );
  AOI21_X1 U143 ( .B1(n807), .B2(n800), .A(n887), .ZN(n188) );
  NAND2_X1 U144 ( .A1(n353), .A2(n592), .ZN(n279) );
  OAI22_X1 U145 ( .A1(n508), .A2(n230), .B1(n509), .B2(n229), .ZN(n507) );
  INV_X1 U146 ( .A(n421), .ZN(n509) );
  OAI22_X1 U147 ( .A1(n207), .A2(n279), .B1(n293), .B2(n206), .ZN(n720) );
  OAI22_X1 U148 ( .A1(n205), .A2(n206), .B1(n207), .B2(n208), .ZN(n204) );
  OAI22_X1 U149 ( .A1(n572), .A2(n468), .B1(n571), .B2(n230), .ZN(n716) );
  NAND2_X1 U150 ( .A1(n338), .A2(n308), .ZN(n306) );
  OAI22_X1 U151 ( .A1(n521), .A2(n208), .B1(n597), .B2(n715), .ZN(n740) );
  OAI22_X1 U152 ( .A1(n571), .A2(n532), .B1(n572), .B2(n533), .ZN(n570) );
  INV_X1 U153 ( .A(n515), .ZN(n458) );
  AND2_X1 U154 ( .A1(n807), .A2(n795), .ZN(n338) );
  NOR2_X1 U155 ( .A1(n478), .A2(n357), .ZN(n548) );
  NAND2_X1 U156 ( .A1(n799), .A2(n810), .ZN(n187) );
  NAND4_X1 U157 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(res[6]) );
  AOI222_X1 U158 ( .A1(N535), .A2(n880), .B1(N635), .B2(n876), .C1(N600), .C2(
        n873), .ZN(n261) );
  AOI222_X1 U159 ( .A1(n225), .A2(n272), .B1(n179), .B2(n273), .C1(n191), .C2(
        n274), .ZN(n263) );
  AOI221_X1 U160 ( .B1(n885), .B2(n275), .C1(N568), .C2(n882), .A(n276), .ZN(
        n262) );
  NAND4_X1 U161 ( .A1(n645), .A2(n646), .A3(n647), .A4(n648), .ZN(res[17]) );
  AOI222_X1 U162 ( .A1(N546), .A2(n881), .B1(N646), .B2(n877), .C1(N611), .C2(
        n875), .ZN(n645) );
  AOI222_X1 U163 ( .A1(n885), .A2(n419), .B1(n515), .B2(n611), .C1(n472), .C2(
        n610), .ZN(n647) );
  AOI221_X1 U164 ( .B1(n191), .B2(n506), .C1(N579), .C2(n882), .A(n656), .ZN(
        n646) );
  NAND4_X1 U165 ( .A1(n766), .A2(n767), .A3(n768), .A4(n769), .ZN(res[10]) );
  AOI222_X1 U166 ( .A1(N539), .A2(n879), .B1(N639), .B2(n878), .C1(N604), .C2(
        n873), .ZN(n766) );
  AOI221_X1 U167 ( .B1(n191), .B2(n275), .C1(n225), .C2(n563), .A(n775), .ZN(
        n768) );
  AOI221_X1 U168 ( .B1(n885), .B2(n483), .C1(N572), .C2(n882), .A(n780), .ZN(
        n767) );
  NAND4_X1 U169 ( .A1(n631), .A2(n632), .A3(n633), .A4(n634), .ZN(res[18]) );
  AOI222_X1 U170 ( .A1(N547), .A2(n881), .B1(N647), .B2(n878), .C1(N612), .C2(
        n875), .ZN(n631) );
  AOI221_X1 U171 ( .B1(n191), .B2(n488), .C1(N580), .C2(n882), .A(n643), .ZN(
        n632) );
  AOI222_X1 U172 ( .A1(n885), .A2(n383), .B1(n515), .B2(n403), .C1(n472), .C2(
        n404), .ZN(n633) );
  NAND4_X1 U173 ( .A1(n312), .A2(n313), .A3(n314), .A4(n315), .ZN(res[3]) );
  AOI222_X1 U174 ( .A1(N532), .A2(n880), .B1(N632), .B2(n877), .C1(N597), .C2(
        n873), .ZN(n312) );
  AOI222_X1 U175 ( .A1(n225), .A2(n254), .B1(n221), .B2(n329), .C1(n179), .C2(
        n330), .ZN(n314) );
  AOI222_X1 U176 ( .A1(N565), .A2(n884), .B1(n193), .B2(n331), .C1(n885), .C2(
        n256), .ZN(n313) );
  NAND4_X1 U177 ( .A1(n238), .A2(n239), .A3(n240), .A4(n241), .ZN(res[7]) );
  AOI222_X1 U178 ( .A1(N536), .A2(n879), .B1(N636), .B2(n876), .C1(N601), .C2(
        n873), .ZN(n238) );
  AOI222_X1 U179 ( .A1(n193), .A2(n254), .B1(n179), .B2(n255), .C1(n191), .C2(
        n256), .ZN(n240) );
  AOI221_X1 U180 ( .B1(n885), .B2(n257), .C1(N569), .C2(n882), .A(n258), .ZN(
        n239) );
  NAND4_X1 U181 ( .A1(n390), .A2(n391), .A3(n392), .A4(n393), .ZN(res[2]) );
  AOI222_X1 U182 ( .A1(N531), .A2(n880), .B1(N631), .B2(n877), .C1(N596), .C2(
        n873), .ZN(n390) );
  AOI222_X1 U183 ( .A1(n225), .A2(n402), .B1(n221), .B2(n403), .C1(n179), .C2(
        n404), .ZN(n392) );
  AOI222_X1 U184 ( .A1(N564), .A2(n884), .B1(n193), .B2(n405), .C1(n885), .C2(
        n274), .ZN(n391) );
  NAND4_X1 U185 ( .A1(n615), .A2(n616), .A3(n617), .A4(n618), .ZN(res[19]) );
  AOI222_X1 U186 ( .A1(N548), .A2(n881), .B1(N648), .B2(n877), .C1(N613), .C2(
        n874), .ZN(n615) );
  AOI222_X1 U187 ( .A1(n885), .A2(n350), .B1(n515), .B2(n329), .C1(n472), .C2(
        n330), .ZN(n617) );
  AOI221_X1 U188 ( .B1(n191), .B2(n629), .C1(N581), .C2(n882), .A(n630), .ZN(
        n616) );
  NAND4_X1 U189 ( .A1(n544), .A2(n545), .A3(n546), .A4(n547), .ZN(res[22]) );
  AOI222_X1 U190 ( .A1(N551), .A2(n880), .B1(N651), .B2(n877), .C1(N616), .C2(
        n874), .ZN(n544) );
  AOI221_X1 U191 ( .B1(n472), .B2(n273), .C1(n885), .C2(n385), .A(n553), .ZN(
        n546) );
  AOI221_X1 U192 ( .B1(n548), .B2(n274), .C1(n549), .C2(n275), .A(n550), .ZN(
        n547) );
  NAND4_X1 U193 ( .A1(n657), .A2(n658), .A3(n659), .A4(n660), .ZN(res[16]) );
  AOI222_X1 U194 ( .A1(N545), .A2(n881), .B1(N645), .B2(n878), .C1(N610), .C2(
        n874), .ZN(n657) );
  AOI222_X1 U195 ( .A1(n191), .A2(n445), .B1(n198), .B2(n224), .C1(n487), .C2(
        n666), .ZN(n659) );
  AOI222_X1 U196 ( .A1(N578), .A2(n884), .B1(n885), .B2(n442), .C1(n667), .C2(
        n592), .ZN(n658) );
  NAND4_X1 U197 ( .A1(n280), .A2(n281), .A3(n282), .A4(n283), .ZN(res[5]) );
  AOI222_X1 U198 ( .A1(N534), .A2(n880), .B1(N634), .B2(n877), .C1(N599), .C2(
        n874), .ZN(n280) );
  AOI221_X1 U199 ( .B1(n221), .B2(n284), .C1(n179), .C2(n285), .A(n286), .ZN(
        n283) );
  AOI221_X1 U200 ( .B1(n885), .B2(n192), .C1(N567), .C2(n882), .A(n292), .ZN(
        n281) );
  NAND4_X1 U201 ( .A1(n704), .A2(n705), .A3(n706), .A4(n707), .ZN(res[13]) );
  AOI221_X1 U202 ( .B1(N607), .B2(n875), .C1(N542), .C2(n879), .A(n725), .ZN(
        n704) );
  AOI221_X1 U203 ( .B1(n191), .B2(n202), .C1(n225), .C2(n500), .A(n716), .ZN(
        n706) );
  AOI221_X1 U204 ( .B1(n200), .B2(n294), .C1(n885), .C2(n506), .A(n720), .ZN(
        n705) );
  NAND4_X1 U205 ( .A1(n686), .A2(n687), .A3(n688), .A4(n689), .ZN(res[14]) );
  AOI221_X1 U206 ( .B1(N608), .B2(n875), .C1(N543), .C2(n879), .A(n702), .ZN(
        n686) );
  AOI221_X1 U207 ( .B1(n198), .B2(n275), .C1(n487), .C2(n274), .A(n697), .ZN(
        n688) );
  AOI221_X1 U208 ( .B1(n225), .B2(n562), .C1(n193), .C2(n563), .A(n700), .ZN(
        n687) );
  NAND2_X1 U209 ( .A1(n796), .A2(n807), .ZN(n362) );
  AOI21_X1 U210 ( .B1(n899), .B2(n246), .A(n892), .ZN(n247) );
  NAND4_X1 U211 ( .A1(n170), .A2(n171), .A3(n172), .A4(n173), .ZN(n164) );
  NOR4_X1 U212 ( .A1(res[30]), .A2(res[2]), .A3(res[29]), .A4(res[28]), .ZN(
        n171) );
  NOR4_X1 U213 ( .A1(res[5]), .A2(res[4]), .A3(res[3]), .A4(res[31]), .ZN(n172) );
  NOR4_X1 U214 ( .A1(res[27]), .A2(res[26]), .A3(res[25]), .A4(res[24]), .ZN(
        n170) );
  NAND2_X1 U215 ( .A1(n799), .A2(n807), .ZN(n434) );
  AOI21_X1 U216 ( .B1(N557), .B2(n879), .A(n389), .ZN(n425) );
  AOI21_X1 U217 ( .B1(N559), .B2(n879), .A(n389), .ZN(n365) );
  NAND4_X1 U218 ( .A1(n745), .A2(n746), .A3(n747), .A4(n748), .ZN(res[11]) );
  AOI22_X1 U219 ( .A1(N573), .A2(n883), .B1(N640), .B2(n876), .ZN(n746) );
  AOI22_X1 U220 ( .A1(N605), .A2(n873), .B1(N540), .B2(n879), .ZN(n745) );
  AOI221_X1 U221 ( .B1(n232), .B2(n254), .C1(n193), .C2(n625), .A(n761), .ZN(
        n747) );
  NAND4_X1 U222 ( .A1(n670), .A2(n671), .A3(n672), .A4(n673), .ZN(res[15]) );
  AOI22_X1 U223 ( .A1(N577), .A2(n883), .B1(N644), .B2(n876), .ZN(n671) );
  AOI22_X1 U224 ( .A1(N609), .A2(n873), .B1(N544), .B2(n879), .ZN(n670) );
  NOR3_X1 U225 ( .A1(n674), .A2(n675), .A3(n676), .ZN(n673) );
  NAND2_X1 U226 ( .A1(n800), .A2(n810), .ZN(n189) );
  OAI21_X1 U227 ( .B1(n551), .B2(n522), .A(n470), .ZN(n550) );
  AOI21_X1 U228 ( .B1(n899), .B2(n552), .A(n892), .ZN(n551) );
  INV_X1 U229 ( .A(n472), .ZN(n463) );
  NAND2_X1 U230 ( .A1(n795), .A2(n810), .ZN(n190) );
  INV_X1 U231 ( .A(n806), .ZN(n796) );
  INV_X1 U232 ( .A(n525), .ZN(n524) );
  AOI22_X1 U233 ( .A1(n442), .A2(n198), .B1(n444), .B2(n191), .ZN(n525) );
  INV_X1 U234 ( .A(n644), .ZN(n643) );
  AOI22_X1 U235 ( .A1(n275), .A2(n487), .B1(n483), .B2(n198), .ZN(n644) );
  AOI221_X1 U236 ( .B1(N763), .B2(n795), .C1(N765), .C2(n796), .A(n797), .ZN(
        n793) );
  INV_X1 U237 ( .A(n798), .ZN(n797) );
  AOI22_X1 U238 ( .A1(N764), .A2(n799), .B1(N762), .B2(n800), .ZN(n798) );
  NAND2_X1 U239 ( .A1(n824), .A2(n799), .ZN(n827) );
  NAND2_X1 U240 ( .A1(n824), .A2(n800), .ZN(n826) );
  AOI21_X1 U241 ( .B1(n804), .B2(n805), .A(n801), .ZN(n803) );
  AOI22_X1 U242 ( .A1(N760), .A2(n799), .B1(N758), .B2(n800), .ZN(n804) );
  AOI22_X1 U243 ( .A1(N759), .A2(n795), .B1(N761), .B2(n796), .ZN(n805) );
  INV_X1 U244 ( .A(n478), .ZN(n452) );
  AND2_X1 U245 ( .A1(n824), .A2(n796), .ZN(n210) );
  AND2_X1 U246 ( .A1(n824), .A2(n795), .ZN(n203) );
  INV_X1 U247 ( .A(n336), .ZN(n335) );
  AOI22_X1 U248 ( .A1(n881), .A2(N560), .B1(n875), .B2(N625), .ZN(n336) );
  INV_X1 U249 ( .A(n726), .ZN(n725) );
  AOI22_X1 U250 ( .A1(N575), .A2(n883), .B1(N642), .B2(n876), .ZN(n726) );
  INV_X1 U251 ( .A(n703), .ZN(n702) );
  AOI22_X1 U252 ( .A1(N576), .A2(n883), .B1(N643), .B2(n876), .ZN(n703) );
  AOI222_X1 U253 ( .A1(n194), .A2(n843), .B1(n500), .B2(n353), .C1(n581), .C2(
        n850), .ZN(n653) );
  AOI222_X1 U254 ( .A1(n272), .A2(n842), .B1(n563), .B2(n853), .C1(n562), .C2(
        n353), .ZN(n640) );
  OAI222_X1 U255 ( .A1(n433), .A2(n461), .B1(n593), .B2(n359), .C1(n521), .C2(
        n357), .ZN(n300) );
  AOI221_X1 U256 ( .B1(n370), .B2(n853), .C1(n562), .C2(n838), .A(n503), .ZN(
        n490) );
  INV_X1 U257 ( .A(n353), .ZN(n461) );
  OAI22_X1 U258 ( .A1(n433), .A2(n357), .B1(n521), .B2(n359), .ZN(n220) );
  OAI221_X1 U259 ( .B1(n521), .B2(n461), .C1(n433), .C2(n639), .A(n811), .ZN(
        n667) );
  AOI22_X1 U260 ( .A1(n844), .A2(n237), .B1(n848), .B2(n226), .ZN(n811) );
  OAI21_X1 U261 ( .B1(n861), .B2(n712), .A(n713), .ZN(n412) );
  NOR2_X1 U262 ( .A1(n712), .A2(n834), .ZN(n346) );
  NOR2_X1 U263 ( .A1(n774), .A2(n834), .ZN(n661) );
  OAI221_X1 U264 ( .B1(n816), .B2(n461), .C1(n744), .C2(n639), .A(n817), .ZN(
        n808) );
  INV_X1 U265 ( .A(n236), .ZN(n816) );
  AOI22_X1 U266 ( .A1(n844), .A2(n818), .B1(n851), .B2(n311), .ZN(n817) );
  NOR2_X1 U267 ( .A1(n624), .A2(n712), .ZN(n503) );
  OAI21_X1 U268 ( .B1(n711), .B2(n712), .A(n713), .ZN(n410) );
  AOI22_X1 U269 ( .A1(n562), .A2(n848), .B1(n563), .B2(n842), .ZN(n557) );
  AOI22_X1 U270 ( .A1(n625), .A2(n838), .B1(n626), .B2(n850), .ZN(n623) );
  AOI22_X1 U271 ( .A1(n581), .A2(n839), .B1(n500), .B2(n849), .ZN(n577) );
  AOI22_X1 U272 ( .A1(n500), .A2(n837), .B1(n412), .B2(n850), .ZN(n182) );
  AOI22_X1 U273 ( .A1(n562), .A2(n840), .B1(n373), .B2(n851), .ZN(n480) );
  NOR2_X1 U274 ( .A1(n834), .A2(n349), .ZN(n380) );
  OAI22_X1 U275 ( .A1(n862), .A2(n381), .B1(n861), .B2(n441), .ZN(n440) );
  OAI22_X1 U276 ( .A1(n862), .A2(n348), .B1(n860), .B2(n381), .ZN(n418) );
  OAI211_X1 U277 ( .C1(n580), .C2(n461), .A(n561), .B(n577), .ZN(n285) );
  OAI211_X1 U278 ( .C1(n540), .C2(n461), .A(n561), .B(n623), .ZN(n330) );
  OAI22_X1 U279 ( .A1(n381), .A2(n872), .B1(n862), .B2(n382), .ZN(n379) );
  OAI22_X1 U280 ( .A1(n872), .A2(n348), .B1(n862), .B2(n349), .ZN(n345) );
  OAI211_X1 U281 ( .C1(n560), .C2(n461), .A(n561), .B(n557), .ZN(n273) );
  AOI21_X1 U282 ( .B1(n353), .B2(n346), .A(n537), .ZN(n253) );
  INV_X1 U283 ( .A(n572), .ZN(n197) );
  OAI21_X1 U284 ( .B1(n556), .B2(n461), .A(n557), .ZN(n266) );
  OAI21_X1 U285 ( .B1(n457), .B2(n624), .A(n623), .ZN(n329) );
  OAI21_X1 U286 ( .B1(n556), .B2(n639), .A(n640), .ZN(n403) );
  OAI21_X1 U287 ( .B1(n560), .B2(n639), .A(n640), .ZN(n404) );
  NAND2_X1 U288 ( .A1(n842), .A2(n308), .ZN(n343) );
  INV_X1 U289 ( .A(n257), .ZN(n462) );
  OAI22_X1 U290 ( .A1(n828), .A2(n826), .B1(n827), .B2(n829), .ZN(N767) );
  NAND2_X1 U291 ( .A1(n830), .A2(n364), .ZN(n829) );
  INV_X1 U292 ( .A(n832), .ZN(n828) );
  XNOR2_X1 U293 ( .A(n712), .B(N625), .ZN(n830) );
  INV_X1 U294 ( .A(n542), .ZN(n356) );
  INV_X1 U295 ( .A(n256), .ZN(n460) );
  INV_X1 U296 ( .A(n451), .ZN(n540) );
  INV_X1 U297 ( .A(n629), .ZN(n358) );
  INV_X1 U298 ( .A(n192), .ZN(n571) );
  INV_X1 U299 ( .A(n736), .ZN(n433) );
  INV_X1 U300 ( .A(n224), .ZN(n519) );
  INV_X1 U301 ( .A(n488), .ZN(n388) );
  INV_X1 U302 ( .A(n202), .ZN(n423) );
  INV_X1 U303 ( .A(n483), .ZN(n387) );
  INV_X1 U304 ( .A(n666), .ZN(n228) );
  INV_X1 U305 ( .A(n402), .ZN(n278) );
  INV_X1 U306 ( .A(n207), .ZN(n581) );
  INV_X1 U307 ( .A(n506), .ZN(n424) );
  INV_X1 U308 ( .A(n445), .ZN(n597) );
  INV_X1 U309 ( .A(n226), .ZN(n593) );
  INV_X1 U310 ( .A(n556), .ZN(n373) );
  INV_X1 U311 ( .A(n194), .ZN(n293) );
  INV_X1 U312 ( .A(n625), .ZN(n260) );
  INV_X1 U313 ( .A(n294), .ZN(n205) );
  INV_X1 U314 ( .A(n383), .ZN(n491) );
  INV_X1 U315 ( .A(n350), .ZN(n469) );
  INV_X1 U316 ( .A(n419), .ZN(n508) );
  INV_X1 U317 ( .A(n272), .ZN(n701) );
  INV_X1 U318 ( .A(n233), .ZN(n744) );
  INV_X1 U319 ( .A(n626), .ZN(n541) );
  INV_X1 U320 ( .A(n502), .ZN(n180) );
  AOI221_X1 U321 ( .B1(n500), .B2(n837), .C1(n410), .C2(n847), .A(n503), .ZN(
        n502) );
  INV_X1 U322 ( .A(n405), .ZN(n277) );
  INV_X1 U323 ( .A(n331), .ZN(n259) );
  INV_X1 U324 ( .A(n560), .ZN(n370) );
  INV_X1 U325 ( .A(n344), .ZN(n326) );
  INV_X1 U326 ( .A(n446), .ZN(n307) );
  INV_X1 U327 ( .A(n242), .ZN(n319) );
  INV_X1 U328 ( .A(n265), .ZN(n397) );
  NOR3_X1 U329 ( .A1(alu_op[3]), .A2(alu_op[4]), .A3(alu_op[2]), .ZN(n807) );
  NOR2_X1 U330 ( .A1(n434), .A2(n694), .ZN(n515) );
  NOR3_X1 U331 ( .A1(alu_op[2]), .A2(alu_op[4]), .A3(n790), .ZN(n810) );
  NOR2_X1 U332 ( .A1(alu_op[0]), .A2(alu_op[1]), .ZN(n800) );
  NOR2_X1 U333 ( .A1(n825), .A2(alu_op[0]), .ZN(n799) );
  AOI222_X1 U334 ( .A1(N629), .A2(n878), .B1(n661), .B2(n885), .C1(N562), .C2(
        n884), .ZN(n785) );
  NOR4_X1 U335 ( .A1(n749), .A2(n750), .A3(n735), .A4(n751), .ZN(n748) );
  NOR3_X1 U336 ( .A1(n183), .A2(b[3]), .A3(n457), .ZN(n751) );
  OAI221_X1 U337 ( .B1(n462), .B2(n229), .C1(n541), .C2(n208), .A(n756), .ZN(
        n749) );
  OAI22_X1 U338 ( .A1(n540), .A2(n693), .B1(n753), .B2(n612), .ZN(n750) );
  AOI221_X1 U339 ( .B1(b[10]), .B2(n770), .C1(n198), .C2(n274), .A(n771), .ZN(
        n769) );
  OAI221_X1 U340 ( .B1(n189), .B2(n613), .C1(a[10]), .C2(n895), .A(n886), .ZN(
        n770) );
  OAI22_X1 U341 ( .A1(n480), .A2(n183), .B1(n772), .B2(n613), .ZN(n771) );
  INV_X1 U342 ( .A(n773), .ZN(n772) );
  AOI221_X1 U343 ( .B1(n549), .B2(n274), .C1(b[18]), .C2(n635), .A(n636), .ZN(
        n634) );
  OAI221_X1 U344 ( .B1(n888), .B2(n594), .C1(a[18]), .C2(n895), .A(n886), .ZN(
        n635) );
  OAI21_X1 U345 ( .B1(n637), .B2(n594), .A(n470), .ZN(n636) );
  INV_X1 U346 ( .A(n638), .ZN(n637) );
  AOI221_X1 U347 ( .B1(n549), .B2(n256), .C1(b[19]), .C2(n619), .A(n620), .ZN(
        n618) );
  OAI221_X1 U348 ( .B1(n888), .B2(n578), .C1(a[19]), .C2(n895), .A(n886), .ZN(
        n619) );
  OAI21_X1 U349 ( .B1(n621), .B2(n578), .A(n470), .ZN(n620) );
  INV_X1 U350 ( .A(n622), .ZN(n621) );
  AOI221_X1 U351 ( .B1(n369), .B2(n451), .C1(n452), .C2(n453), .A(n454), .ZN(
        n450) );
  OAI222_X1 U352 ( .A1(n460), .A2(n461), .B1(n356), .B2(n359), .C1(n462), .C2(
        n357), .ZN(n453) );
  OAI21_X1 U353 ( .B1(n455), .B2(n381), .A(n456), .ZN(n454) );
  OR3_X1 U354 ( .A1(n457), .A2(b[3]), .A3(n458), .ZN(n456) );
  AOI221_X1 U355 ( .B1(n200), .B2(n265), .C1(n221), .C2(n266), .A(n267), .ZN(
        n264) );
  OAI22_X1 U356 ( .A1(n268), .A2(n269), .B1(n270), .B2(n271), .ZN(n267) );
  AOI221_X1 U357 ( .B1(n897), .B2(n271), .C1(a[6]), .C2(n889), .A(n887), .ZN(
        n268) );
  AOI21_X1 U358 ( .B1(n898), .B2(n269), .A(n892), .ZN(n270) );
  AOI221_X1 U359 ( .B1(n682), .B2(n373), .C1(b[14]), .C2(n690), .A(n691), .ZN(
        n689) );
  OAI221_X1 U360 ( .B1(n189), .B2(n668), .C1(a[14]), .C2(n895), .A(n886), .ZN(
        n690) );
  OAI221_X1 U361 ( .B1(n692), .B2(n668), .C1(n560), .C2(n693), .A(n695), .ZN(
        n691) );
  INV_X1 U362 ( .A(n696), .ZN(n692) );
  AOI221_X1 U363 ( .B1(n200), .B2(n242), .C1(n221), .C2(n243), .A(n244), .ZN(
        n241) );
  INV_X1 U364 ( .A(n253), .ZN(n243) );
  OAI22_X1 U365 ( .A1(n245), .A2(n246), .B1(n247), .B2(n248), .ZN(n244) );
  AOI221_X1 U366 ( .B1(n897), .B2(n248), .C1(a[7]), .C2(n889), .A(n887), .ZN(
        n245) );
  AOI221_X1 U367 ( .B1(a[2]), .B2(n394), .C1(b[2]), .C2(n395), .A(n396), .ZN(
        n393) );
  OAI221_X1 U368 ( .B1(n888), .B2(n401), .C1(a[2]), .C2(n894), .A(n886), .ZN(
        n395) );
  OAI21_X1 U369 ( .B1(b[2]), .B2(n893), .A(n891), .ZN(n394) );
  OAI22_X1 U370 ( .A1(n397), .A2(n206), .B1(n398), .B2(n321), .ZN(n396) );
  AOI221_X1 U371 ( .B1(a[3]), .B2(n316), .C1(b[3]), .C2(n317), .A(n318), .ZN(
        n315) );
  OAI221_X1 U372 ( .B1(n888), .B2(n328), .C1(a[3]), .C2(n894), .A(n886), .ZN(
        n317) );
  OAI21_X1 U373 ( .B1(b[3]), .B2(n893), .A(n891), .ZN(n316) );
  OAI22_X1 U374 ( .A1(n319), .A2(n206), .B1(n320), .B2(n321), .ZN(n318) );
  AOI221_X1 U375 ( .B1(n731), .B2(n446), .C1(a[12]), .C2(n732), .A(n733), .ZN(
        n730) );
  NOR2_X1 U376 ( .A1(n624), .A2(n306), .ZN(n731) );
  OAI21_X1 U377 ( .B1(b[12]), .B2(n893), .A(n890), .ZN(n732) );
  NAND2_X1 U378 ( .A1(n734), .A2(n695), .ZN(n733) );
  AOI221_X1 U379 ( .B1(n682), .B2(n412), .C1(b[13]), .C2(n708), .A(n709), .ZN(
        n707) );
  OAI221_X1 U380 ( .B1(n189), .B2(n678), .C1(a[13]), .C2(n895), .A(n886), .ZN(
        n708) );
  OAI221_X1 U381 ( .B1(n710), .B2(n678), .C1(n580), .C2(n693), .A(n695), .ZN(
        n709) );
  INV_X1 U382 ( .A(n714), .ZN(n710) );
  AOI221_X1 U383 ( .B1(n549), .B2(n197), .C1(b[17]), .C2(n649), .A(n650), .ZN(
        n648) );
  OAI221_X1 U384 ( .B1(n888), .B2(n627), .C1(a[17]), .C2(n895), .A(n886), .ZN(
        n649) );
  OAI21_X1 U385 ( .B1(n651), .B2(n627), .A(n470), .ZN(n650) );
  INV_X1 U386 ( .A(n652), .ZN(n651) );
  AOI221_X1 U387 ( .B1(n549), .B2(n661), .C1(b[16]), .C2(n662), .A(n663), .ZN(
        n660) );
  OAI221_X1 U388 ( .B1(n888), .B2(n641), .C1(a[16]), .C2(n895), .A(n886), .ZN(
        n662) );
  OAI21_X1 U389 ( .B1(n664), .B2(n641), .A(n470), .ZN(n663) );
  INV_X1 U390 ( .A(n665), .ZN(n664) );
  AOI211_X1 U391 ( .C1(n587), .C2(n452), .A(n588), .B(n309), .ZN(n586) );
  NOR2_X1 U392 ( .A1(b[3]), .A2(n307), .ZN(n587) );
  OAI22_X1 U393 ( .A1(n463), .A2(n561), .B1(n589), .B2(n558), .ZN(n588) );
  INV_X1 U394 ( .A(n590), .ZN(n589) );
  OAI221_X1 U395 ( .B1(n888), .B2(n558), .C1(a[20]), .C2(n894), .A(n886), .ZN(
        n591) );
  OAI221_X1 U396 ( .B1(n888), .B2(n485), .C1(a[24]), .C2(n894), .A(n886), .ZN(
        n520) );
  OAI221_X1 U397 ( .B1(n465), .B2(n189), .C1(a[25]), .C2(n894), .A(n886), .ZN(
        n501) );
  OAI221_X1 U398 ( .B1(n441), .B2(n189), .C1(a[26]), .C2(n894), .A(n886), .ZN(
        n484) );
  OAI221_X1 U399 ( .B1(n888), .B2(n774), .C1(a[0]), .C2(n893), .A(n886), .ZN(
        n809) );
  OAI221_X1 U400 ( .B1(n888), .B2(n223), .C1(a[8]), .C2(n894), .A(n886), .ZN(
        n216) );
  OAI221_X1 U401 ( .B1(n348), .B2(n189), .C1(a[28]), .C2(n894), .A(n886), .ZN(
        n429) );
  OAI22_X1 U402 ( .A1(n605), .A2(n206), .B1(n606), .B2(n321), .ZN(n604) );
  INV_X1 U403 ( .A(n291), .ZN(n605) );
  AOI221_X1 U404 ( .B1(a[4]), .B2(n322), .C1(a[1]), .C2(n867), .A(n607), .ZN(
        n606) );
  OAI22_X1 U405 ( .A1(n862), .A2(n401), .B1(n860), .B2(n328), .ZN(n607) );
  OAI22_X1 U406 ( .A1(n182), .A2(n183), .B1(n184), .B2(n185), .ZN(n181) );
  INV_X1 U407 ( .A(n186), .ZN(n184) );
  OAI21_X1 U408 ( .B1(n894), .B2(b[9]), .A(n891), .ZN(n186) );
  NAND2_X1 U409 ( .A1(n338), .A2(n694), .ZN(n478) );
  AOI22_X1 U410 ( .A1(b[11]), .A2(n757), .B1(n198), .B2(n256), .ZN(n756) );
  OAI221_X1 U411 ( .B1(n189), .B2(n612), .C1(a[11]), .C2(n895), .A(n886), .ZN(
        n757) );
  NAND4_X1 U412 ( .A1(n583), .A2(n584), .A3(n585), .A4(n586), .ZN(res[20]) );
  AOI222_X1 U413 ( .A1(N549), .A2(n880), .B1(N649), .B2(n877), .C1(N614), .C2(
        n874), .ZN(n583) );
  AOI222_X1 U414 ( .A1(n885), .A2(n444), .B1(b[20]), .B2(n591), .C1(n592), 
        .C2(n300), .ZN(n585) );
  AOI221_X1 U415 ( .B1(n191), .B2(n442), .C1(N582), .C2(n883), .A(n596), .ZN(
        n584) );
  NAND4_X1 U416 ( .A1(n510), .A2(n511), .A3(n512), .A4(n513), .ZN(res[24]) );
  AOI222_X1 U417 ( .A1(N553), .A2(n880), .B1(N653), .B2(n877), .C1(N618), .C2(
        n874), .ZN(n510) );
  AOI222_X1 U418 ( .A1(n885), .A2(n443), .B1(b[24]), .B2(n520), .C1(n472), 
        .C2(n217), .ZN(n512) );
  AOI221_X1 U419 ( .B1(n487), .B2(n445), .C1(N586), .C2(n883), .A(n524), .ZN(
        n511) );
  NAND4_X1 U420 ( .A1(n565), .A2(n566), .A3(n567), .A4(n568), .ZN(res[21]) );
  AOI222_X1 U421 ( .A1(N550), .A2(n880), .B1(N650), .B2(n877), .C1(N615), .C2(
        n874), .ZN(n565) );
  AOI211_X1 U422 ( .C1(a[21]), .C2(n569), .A(n570), .B(n309), .ZN(n568) );
  AOI221_X1 U423 ( .B1(n472), .B2(n285), .C1(n885), .C2(n421), .A(n573), .ZN(
        n567) );
  NAND4_X1 U424 ( .A1(n492), .A2(n493), .A3(n494), .A4(n495), .ZN(res[25]) );
  AOI222_X1 U425 ( .A1(N554), .A2(n880), .B1(N654), .B2(n877), .C1(N619), .C2(
        n874), .ZN(n492) );
  AOI222_X1 U426 ( .A1(n885), .A2(n420), .B1(b[25]), .B2(n501), .C1(n472), 
        .C2(n180), .ZN(n494) );
  AOI221_X1 U427 ( .B1(n487), .B2(n506), .C1(N587), .C2(n882), .A(n507), .ZN(
        n493) );
  NAND4_X1 U428 ( .A1(n295), .A2(n296), .A3(n297), .A4(n298), .ZN(res[4]) );
  AOI222_X1 U429 ( .A1(N533), .A2(n880), .B1(N633), .B2(n876), .C1(N598), .C2(
        n873), .ZN(n295) );
  AOI221_X1 U430 ( .B1(n299), .B2(n300), .C1(n694), .C2(n301), .A(n302), .ZN(
        n298) );
  AOI222_X1 U431 ( .A1(N566), .A2(n884), .B1(n200), .B2(n311), .C1(n232), .C2(
        n236), .ZN(n296) );
  NAND4_X1 U432 ( .A1(n212), .A2(n213), .A3(n214), .A4(n215), .ZN(res[8]) );
  AOI222_X1 U433 ( .A1(N537), .A2(n879), .B1(N637), .B2(n876), .C1(N602), .C2(
        n873), .ZN(n212) );
  AOI221_X1 U434 ( .B1(b[8]), .B2(n216), .C1(n179), .C2(n217), .A(n218), .ZN(
        n215) );
  AOI221_X1 U435 ( .B1(n885), .B2(n224), .C1(n225), .C2(n226), .A(n227), .ZN(
        n214) );
  NAND4_X1 U436 ( .A1(n473), .A2(n474), .A3(n475), .A4(n476), .ZN(res[26]) );
  AOI222_X1 U437 ( .A1(N555), .A2(n880), .B1(N655), .B2(n877), .C1(N620), .C2(
        n874), .ZN(n473) );
  AOI222_X1 U438 ( .A1(n191), .A2(n385), .B1(b[26]), .B2(n484), .C1(n885), 
        .C2(n384), .ZN(n475) );
  AOI221_X1 U439 ( .B1(n487), .B2(n488), .C1(N588), .C2(n882), .A(n489), .ZN(
        n474) );
  NAND4_X1 U440 ( .A1(n598), .A2(n599), .A3(n600), .A4(n601), .ZN(res[1]) );
  AOI222_X1 U441 ( .A1(N530), .A2(n881), .B1(N630), .B2(n878), .C1(N595), .C2(
        n874), .ZN(n598) );
  AOI222_X1 U442 ( .A1(n179), .A2(n610), .B1(n193), .B2(n199), .C1(n221), .C2(
        n611), .ZN(n600) );
  AOI221_X1 U443 ( .B1(a[1]), .B2(n602), .C1(b[1]), .C2(n603), .A(n604), .ZN(
        n601) );
  NAND4_X1 U444 ( .A1(n727), .A2(n728), .A3(n729), .A4(n730), .ZN(res[12]) );
  AOI222_X1 U445 ( .A1(N541), .A2(n881), .B1(N641), .B2(n878), .C1(N606), .C2(
        n874), .ZN(n727) );
  AOI221_X1 U446 ( .B1(b[12]), .B2(n739), .C1(n191), .C2(n224), .A(n740), .ZN(
        n729) );
  AOI221_X1 U447 ( .B1(n232), .B2(n237), .C1(N574), .C2(n882), .A(n743), .ZN(
        n728) );
  NAND4_X1 U448 ( .A1(n174), .A2(n175), .A3(n176), .A4(n177), .ZN(res[9]) );
  AOI222_X1 U449 ( .A1(N538), .A2(n880), .B1(N638), .B2(n876), .C1(N603), .C2(
        n873), .ZN(n174) );
  AOI221_X1 U450 ( .B1(b[9]), .B2(n178), .C1(n179), .C2(n180), .A(n181), .ZN(
        n177) );
  AOI221_X1 U451 ( .B1(n885), .B2(n202), .C1(N571), .C2(n882), .A(n204), .ZN(
        n175) );
  NAND4_X1 U452 ( .A1(n526), .A2(n527), .A3(n528), .A4(n529), .ZN(res[23]) );
  AOI222_X1 U453 ( .A1(N552), .A2(n880), .B1(N652), .B2(n877), .C1(N617), .C2(
        n874), .ZN(n526) );
  AOI221_X1 U454 ( .B1(n472), .B2(n255), .C1(n885), .C2(n354), .A(n534), .ZN(
        n528) );
  AOI211_X1 U455 ( .C1(a[23]), .C2(n530), .A(n531), .B(n309), .ZN(n529) );
  NAND2_X1 U456 ( .A1(n470), .A2(n471), .ZN(n389) );
  OAI211_X1 U457 ( .C1(n834), .C2(n361), .A(n362), .B(n363), .ZN(n337) );
  AOI21_X1 U458 ( .B1(b[31]), .B2(n889), .A(n892), .ZN(n363) );
  NAND4_X1 U459 ( .A1(n447), .A2(n448), .A3(n449), .A4(n450), .ZN(res[27]) );
  AOI222_X1 U460 ( .A1(n191), .A2(n354), .B1(b[27]), .B2(n464), .C1(n885), 
        .C2(n352), .ZN(n449) );
  AOI221_X1 U461 ( .B1(N589), .B2(n884), .C1(N656), .C2(n876), .A(n467), .ZN(
        n448) );
  AOI221_X1 U462 ( .B1(N621), .B2(n875), .C1(N556), .C2(n879), .A(n389), .ZN(
        n447) );
  NAND4_X1 U463 ( .A1(n784), .A2(n785), .A3(n786), .A4(n787), .ZN(res[0]) );
  AOI22_X1 U464 ( .A1(N594), .A2(n873), .B1(N529), .B2(n879), .ZN(n784) );
  AOI222_X1 U465 ( .A1(n808), .A2(n592), .B1(n667), .B2(n299), .C1(b[0]), .C2(
        n809), .ZN(n786) );
  AOI21_X1 U466 ( .B1(a[0]), .B2(n788), .A(n789), .ZN(n787) );
  NAND4_X1 U467 ( .A1(n406), .A2(n407), .A3(n408), .A4(n409), .ZN(res[29]) );
  AOI222_X1 U468 ( .A1(N623), .A2(n875), .B1(N591), .B2(n883), .C1(N658), .C2(
        n878), .ZN(n407) );
  AOI22_X1 U469 ( .A1(b[29]), .A2(n413), .B1(n338), .B2(n414), .ZN(n408) );
  AOI21_X1 U470 ( .B1(N558), .B2(n879), .A(n389), .ZN(n406) );
  OAI22_X1 U471 ( .A1(n287), .A2(n288), .B1(n289), .B2(n290), .ZN(n286) );
  AOI221_X1 U472 ( .B1(n897), .B2(n290), .C1(a[5]), .C2(n889), .A(n887), .ZN(
        n287) );
  AOI21_X1 U473 ( .B1(n899), .B2(n288), .A(n892), .ZN(n289) );
  INV_X1 U474 ( .A(b[5]), .ZN(n288) );
  OAI21_X1 U475 ( .B1(n303), .B2(n304), .A(n305), .ZN(n302) );
  OR3_X1 U476 ( .A1(n306), .A2(b[3]), .A3(n307), .ZN(n305) );
  AOI21_X1 U477 ( .B1(n898), .B2(n308), .A(n892), .ZN(n303) );
  NAND4_X1 U478 ( .A1(n365), .A2(n366), .A3(n367), .A4(n368), .ZN(res[30]) );
  AOI222_X1 U479 ( .A1(N624), .A2(n875), .B1(N592), .B2(n883), .C1(N659), .C2(
        n878), .ZN(n366) );
  AOI22_X1 U480 ( .A1(b[30]), .A2(n374), .B1(n338), .B2(n375), .ZN(n367) );
  AOI222_X1 U481 ( .A1(n369), .A2(n370), .B1(a[30]), .B2(n371), .C1(n372), 
        .C2(n373), .ZN(n368) );
  AOI22_X1 U482 ( .A1(n887), .A2(b[31]), .B1(n898), .B2(n364), .ZN(n332) );
  AOI221_X1 U483 ( .B1(N593), .B2(n884), .C1(N660), .C2(n876), .A(n335), .ZN(
        n334) );
  AOI22_X1 U484 ( .A1(a[31]), .A2(n337), .B1(n338), .B2(n339), .ZN(n333) );
  AND2_X1 U485 ( .A1(alu_op[0]), .A2(n825), .ZN(n795) );
  OAI21_X1 U486 ( .B1(n895), .B2(b[24]), .A(n891), .ZN(n518) );
  OAI21_X1 U487 ( .B1(n896), .B2(b[10]), .A(n890), .ZN(n773) );
  OAI21_X1 U488 ( .B1(n896), .B2(b[13]), .A(n890), .ZN(n714) );
  OAI21_X1 U489 ( .B1(n896), .B2(b[14]), .A(n890), .ZN(n696) );
  OAI21_X1 U490 ( .B1(n896), .B2(b[15]), .A(n890), .ZN(n684) );
  OAI21_X1 U491 ( .B1(n896), .B2(b[16]), .A(n890), .ZN(n665) );
  OAI21_X1 U492 ( .B1(n896), .B2(b[17]), .A(n890), .ZN(n652) );
  OAI21_X1 U493 ( .B1(n896), .B2(b[18]), .A(n890), .ZN(n638) );
  OAI21_X1 U494 ( .B1(n896), .B2(b[19]), .A(n890), .ZN(n622) );
  OAI21_X1 U495 ( .B1(n896), .B2(b[20]), .A(n891), .ZN(n590) );
  OAI21_X1 U496 ( .B1(n895), .B2(b[25]), .A(n891), .ZN(n499) );
  OAI21_X1 U497 ( .B1(n896), .B2(b[26]), .A(n891), .ZN(n482) );
  OAI21_X1 U498 ( .B1(b[28]), .B2(n893), .A(n891), .ZN(n430) );
  OAI21_X1 U499 ( .B1(b[0]), .B2(n893), .A(n890), .ZN(n788) );
  OAI21_X1 U500 ( .B1(b[21]), .B2(n893), .A(n891), .ZN(n569) );
  OAI21_X1 U501 ( .B1(b[23]), .B2(n893), .A(n891), .ZN(n530) );
  OAI21_X1 U502 ( .B1(b[30]), .B2(n893), .A(n891), .ZN(n371) );
  AOI222_X1 U503 ( .A1(n369), .A2(n410), .B1(a[29]), .B2(n411), .C1(n372), 
        .C2(n412), .ZN(n409) );
  OAI21_X1 U504 ( .B1(b[29]), .B2(n893), .A(n891), .ZN(n411) );
  OAI21_X1 U505 ( .B1(b[1]), .B2(n893), .A(n890), .ZN(n602) );
  NAND4_X1 U506 ( .A1(n425), .A2(n426), .A3(n427), .A4(n428), .ZN(res[28]) );
  AOI22_X1 U507 ( .A1(n338), .A2(n435), .B1(N590), .B2(n883), .ZN(n427) );
  AOI22_X1 U508 ( .A1(N657), .A2(n876), .B1(N622), .B2(n873), .ZN(n426) );
  AOI221_X1 U509 ( .B1(b[28]), .B2(n429), .C1(a[28]), .C2(n430), .A(n431), 
        .ZN(n428) );
  INV_X1 U510 ( .A(alu_op[3]), .ZN(n790) );
  NAND2_X1 U511 ( .A1(alu_op[1]), .A2(alu_op[0]), .ZN(n806) );
  INV_X1 U512 ( .A(alu_op[1]), .ZN(n825) );
  INV_X1 U513 ( .A(n477), .ZN(n476) );
  OAI221_X1 U514 ( .B1(n478), .B2(n479), .C1(n458), .C2(n480), .A(n481), .ZN(
        n477) );
  AOI222_X1 U515 ( .A1(n274), .A2(n353), .B1(n483), .B2(n838), .C1(n275), .C2(
        n851), .ZN(n479) );
  AOI21_X1 U516 ( .B1(n482), .B2(a[26]), .A(n309), .ZN(n481) );
  INV_X1 U517 ( .A(n496), .ZN(n495) );
  OAI221_X1 U518 ( .B1(n478), .B2(n497), .C1(n458), .C2(n182), .A(n498), .ZN(
        n496) );
  AOI222_X1 U519 ( .A1(n197), .A2(n353), .B1(n192), .B2(n852), .C1(n202), .C2(
        n840), .ZN(n497) );
  AOI21_X1 U520 ( .B1(n499), .B2(a[25]), .A(n309), .ZN(n498) );
  INV_X1 U521 ( .A(n219), .ZN(n218) );
  AOI22_X1 U522 ( .A1(n220), .A2(n221), .B1(n222), .B2(a[8]), .ZN(n219) );
  OAI21_X1 U523 ( .B1(n896), .B2(b[8]), .A(n891), .ZN(n222) );
  INV_X1 U524 ( .A(n574), .ZN(n573) );
  AOI22_X1 U525 ( .A1(n284), .A2(n515), .B1(n575), .B2(b[21]), .ZN(n574) );
  OAI221_X1 U526 ( .B1(n893), .B2(a[21]), .C1(n538), .C2(n189), .A(n886), .ZN(
        n575) );
  INV_X1 U527 ( .A(n754), .ZN(n753) );
  OAI21_X1 U528 ( .B1(n896), .B2(b[11]), .A(n890), .ZN(n754) );
  INV_X1 U529 ( .A(n459), .ZN(n455) );
  OAI21_X1 U530 ( .B1(n896), .B2(b[27]), .A(n891), .ZN(n459) );
  OAI211_X1 U531 ( .C1(n680), .C2(n654), .A(n470), .B(n681), .ZN(n674) );
  AOI22_X1 U532 ( .A1(n682), .A2(n346), .B1(b[15]), .B2(n683), .ZN(n681) );
  INV_X1 U533 ( .A(n684), .ZN(n680) );
  OAI221_X1 U534 ( .B1(n189), .B2(n654), .C1(a[15]), .C2(n895), .A(n886), .ZN(
        n683) );
  NOR2_X1 U535 ( .A1(n164), .A2(n165), .ZN(zero) );
  NAND4_X1 U536 ( .A1(n166), .A2(n167), .A3(n168), .A4(n169), .ZN(n165) );
  INV_X1 U537 ( .A(alu_op[4]), .ZN(n794) );
  NAND2_X1 U538 ( .A1(n801), .A2(n790), .ZN(n792) );
  AOI21_X1 U539 ( .B1(n802), .B2(N757), .A(n803), .ZN(n791) );
  NOR3_X1 U540 ( .A1(alu_op[3]), .A2(alu_op[4]), .A3(n801), .ZN(n824) );
  OAI221_X1 U541 ( .B1(n888), .B2(n609), .C1(a[1]), .C2(n895), .A(n886), .ZN(
        n603) );
  OAI221_X1 U542 ( .B1(n888), .B2(n304), .C1(a[4]), .C2(n894), .A(n886), .ZN(
        n301) );
  OAI221_X1 U543 ( .B1(n382), .B2(n189), .C1(a[29]), .C2(n894), .A(n886), .ZN(
        n413) );
  OAI221_X1 U544 ( .B1(n349), .B2(n189), .C1(a[30]), .C2(n894), .A(n886), .ZN(
        n374) );
  OAI221_X1 U545 ( .B1(n381), .B2(n189), .C1(a[27]), .C2(n894), .A(n886), .ZN(
        n464) );
  OAI221_X1 U546 ( .B1(n189), .B2(n698), .C1(a[12]), .C2(n895), .A(n886), .ZN(
        n739) );
  OAI221_X1 U547 ( .B1(n185), .B2(n888), .C1(a[9]), .C2(n894), .A(n886), .ZN(
        n178) );
  OAI22_X1 U548 ( .A1(n554), .A2(n458), .B1(n555), .B2(n552), .ZN(n553) );
  INV_X1 U549 ( .A(n266), .ZN(n554) );
  AOI221_X1 U550 ( .B1(n898), .B2(n522), .C1(a[22]), .C2(n889), .A(n887), .ZN(
        n555) );
  OAI22_X1 U551 ( .A1(n253), .A2(n458), .B1(n535), .B2(n536), .ZN(n534) );
  INV_X1 U552 ( .A(b[23]), .ZN(n536) );
  AOI221_X1 U553 ( .B1(n899), .B2(n504), .C1(a[23]), .C2(n889), .A(n887), .ZN(
        n535) );
  NOR2_X1 U554 ( .A1(alu_op[2]), .A2(n806), .ZN(n802) );
  INV_X1 U555 ( .A(alu_op[2]), .ZN(n801) );
  AOI22_X1 U556 ( .A1(a[3]), .A2(n322), .B1(a[6]), .B2(n867), .ZN(n779) );
  OAI22_X1 U557 ( .A1(n872), .A2(n381), .B1(n485), .B2(n834), .ZN(n815) );
  OAI221_X1 U558 ( .B1(n859), .B2(n609), .C1(n863), .C2(n401), .A(n758), .ZN(
        n256) );
  AOI22_X1 U559 ( .A1(a[0]), .A2(n871), .B1(a[3]), .B2(n866), .ZN(n758) );
  OAI221_X1 U560 ( .B1(n859), .B2(n271), .C1(n863), .C2(n248), .A(n742), .ZN(
        n224) );
  AOI22_X1 U561 ( .A1(a[5]), .A2(n871), .B1(a[8]), .B2(n866), .ZN(n742) );
  OAI221_X1 U562 ( .B1(n858), .B2(n381), .C1(n862), .C2(n441), .A(n718), .ZN(
        n500) );
  AOI22_X1 U563 ( .A1(a[28]), .A2(n870), .B1(a[25]), .B2(n866), .ZN(n718) );
  INV_X1 U564 ( .A(N560), .ZN(n833) );
  OAI221_X1 U565 ( .B1(n858), .B2(n328), .C1(n864), .C2(n304), .A(n717), .ZN(
        n192) );
  AOI22_X1 U566 ( .A1(a[2]), .A2(n870), .B1(a[5]), .B2(n867), .ZN(n717) );
  OAI221_X1 U568 ( .B1(n858), .B2(n248), .C1(n863), .C2(n223), .A(n719), .ZN(
        n202) );
  AOI22_X1 U569 ( .A1(a[6]), .A2(n870), .B1(n868), .B2(a[9]), .ZN(n719) );
  OAI221_X1 U570 ( .B1(n859), .B2(n348), .C1(n864), .C2(n381), .A(n782), .ZN(
        n562) );
  AOI22_X1 U571 ( .A1(n869), .A2(a[29]), .B1(a[26]), .B2(n867), .ZN(n782) );
  OAI221_X1 U572 ( .B1(n860), .B2(n223), .C1(n185), .C2(n862), .A(n783), .ZN(
        n483) );
  AOI22_X1 U573 ( .A1(a[7]), .A2(n322), .B1(a[10]), .B2(n867), .ZN(n783) );
  AOI221_X1 U574 ( .B1(n344), .B2(a[23]), .C1(n865), .C2(a[22]), .A(n722), 
        .ZN(n207) );
  OAI22_X1 U575 ( .A1(n485), .A2(n872), .B1(n538), .B2(n834), .ZN(n722) );
  NOR2_X2 U576 ( .A1(n624), .A2(b[2]), .ZN(n353) );
  OAI221_X1 U577 ( .B1(n859), .B2(n627), .C1(n863), .C2(n641), .A(n765), .ZN(
        n254) );
  AOI22_X1 U578 ( .A1(a[18]), .A2(n871), .B1(a[15]), .B2(n867), .ZN(n765) );
  OAI221_X1 U579 ( .B1(n858), .B2(n612), .C1(n325), .C2(n698), .A(n723), .ZN(
        n506) );
  AOI22_X1 U580 ( .A1(a[10]), .A2(n870), .B1(a[13]), .B2(n866), .ZN(n723) );
  OAI221_X1 U581 ( .B1(n860), .B2(n485), .C1(n862), .C2(n504), .A(n778), .ZN(
        n563) );
  AOI22_X1 U582 ( .A1(a[25]), .A2(n871), .B1(a[22]), .B2(n867), .ZN(n778) );
  OAI221_X1 U583 ( .B1(n860), .B2(n594), .C1(n325), .C2(n627), .A(n813), .ZN(
        n237) );
  AOI22_X1 U584 ( .A1(a[19]), .A2(n322), .B1(a[16]), .B2(n868), .ZN(n813) );
  OAI221_X1 U585 ( .B1(n858), .B2(n668), .C1(n864), .C2(n654), .A(n669), .ZN(
        n442) );
  AOI22_X1 U586 ( .A1(a[13]), .A2(n870), .B1(a[16]), .B2(n868), .ZN(n669) );
  OAI221_X1 U587 ( .B1(n859), .B2(n613), .C1(n863), .C2(n612), .A(n741), .ZN(
        n445) );
  AOI22_X1 U588 ( .A1(n871), .A2(a[9]), .B1(a[12]), .B2(n866), .ZN(n741) );
  NOR2_X1 U589 ( .A1(n711), .A2(b[0]), .ZN(n344) );
  OAI221_X1 U590 ( .B1(n860), .B2(n522), .C1(n864), .C2(n538), .A(n812), .ZN(
        n226) );
  AOI22_X1 U591 ( .A1(a[23]), .A2(n322), .B1(a[20]), .B2(n867), .ZN(n812) );
  OAI221_X1 U592 ( .B1(n859), .B2(n578), .C1(n864), .C2(n558), .A(n579), .ZN(
        n421) );
  AOI22_X1 U593 ( .A1(a[18]), .A2(n870), .B1(a[21]), .B2(n866), .ZN(n579) );
  OAI221_X1 U594 ( .B1(n857), .B2(n558), .C1(n864), .C2(n538), .A(n559), .ZN(
        n385) );
  AOI22_X1 U595 ( .A1(a[19]), .A2(n869), .B1(a[22]), .B2(n868), .ZN(n559) );
  OAI221_X1 U596 ( .B1(n857), .B2(n538), .C1(n864), .C2(n522), .A(n539), .ZN(
        n354) );
  AOI22_X1 U597 ( .A1(a[20]), .A2(n869), .B1(a[23]), .B2(n866), .ZN(n539) );
  OAI221_X1 U598 ( .B1(n858), .B2(n578), .C1(n325), .C2(n594), .A(n721), .ZN(
        n194) );
  AOI22_X1 U599 ( .A1(a[20]), .A2(n870), .B1(a[17]), .B2(n866), .ZN(n721) );
  OAI221_X1 U600 ( .B1(n859), .B2(n538), .C1(n863), .C2(n558), .A(n764), .ZN(
        n625) );
  AOI22_X1 U601 ( .A1(a[22]), .A2(n871), .B1(a[19]), .B2(n867), .ZN(n764) );
  OAI221_X1 U602 ( .B1(n859), .B2(n290), .C1(n863), .C2(n271), .A(n760), .ZN(
        n257) );
  AOI22_X1 U603 ( .A1(a[4]), .A2(n871), .B1(a[7]), .B2(n866), .ZN(n760) );
  OAI221_X1 U604 ( .B1(n382), .B2(n861), .C1(n863), .C2(n348), .A(n755), .ZN(
        n451) );
  AOI22_X1 U605 ( .A1(n869), .A2(a[30]), .B1(a[27]), .B2(n866), .ZN(n755) );
  OAI221_X1 U606 ( .B1(n858), .B2(n654), .C1(n325), .C2(n668), .A(n724), .ZN(
        n294) );
  AOI22_X1 U607 ( .A1(a[16]), .A2(n870), .B1(a[13]), .B2(n866), .ZN(n724) );
  OAI221_X1 U608 ( .B1(n857), .B2(n613), .C1(n185), .C2(n862), .A(n822), .ZN(
        n236) );
  AOI22_X1 U609 ( .A1(a[11]), .A2(n869), .B1(a[8]), .B2(n868), .ZN(n822) );
  OAI221_X1 U610 ( .B1(n857), .B2(n612), .C1(n325), .C2(n613), .A(n614), .ZN(
        n199) );
  AOI22_X1 U611 ( .A1(a[12]), .A2(n869), .B1(n868), .B2(a[9]), .ZN(n614) );
  OAI221_X1 U612 ( .B1(n858), .B2(n654), .C1(n325), .C2(n641), .A(n655), .ZN(
        n419) );
  AOI22_X1 U613 ( .A1(a[14]), .A2(n870), .B1(a[17]), .B2(n866), .ZN(n655) );
  OAI221_X1 U614 ( .B1(n858), .B2(n641), .C1(n325), .C2(n627), .A(n642), .ZN(
        n383) );
  AOI22_X1 U615 ( .A1(a[15]), .A2(n870), .B1(a[18]), .B2(n867), .ZN(n642) );
  OAI221_X1 U616 ( .B1(n857), .B2(n627), .C1(n325), .C2(n594), .A(n628), .ZN(
        n350) );
  AOI22_X1 U617 ( .A1(a[16]), .A2(n869), .B1(a[19]), .B2(n868), .ZN(n628) );
  OAI221_X1 U618 ( .B1(n859), .B2(n558), .C1(n863), .C2(n578), .A(n776), .ZN(
        n272) );
  AOI22_X1 U619 ( .A1(a[21]), .A2(n871), .B1(a[18]), .B2(n867), .ZN(n776) );
  OAI221_X1 U620 ( .B1(n860), .B2(n668), .C1(n325), .C2(n678), .A(n821), .ZN(
        n233) );
  AOI22_X1 U621 ( .A1(a[15]), .A2(n871), .B1(a[12]), .B2(n867), .ZN(n821) );
  OAI221_X1 U622 ( .B1(n858), .B2(n698), .C1(n325), .C2(n678), .A(n699), .ZN(
        n488) );
  AOI22_X1 U623 ( .A1(a[11]), .A2(n870), .B1(a[14]), .B2(n868), .ZN(n699) );
  OAI221_X1 U624 ( .B1(n857), .B2(n594), .C1(n864), .C2(n578), .A(n595), .ZN(
        n444) );
  AOI22_X1 U625 ( .A1(a[17]), .A2(n869), .B1(a[20]), .B2(n868), .ZN(n595) );
  OAI221_X1 U626 ( .B1(n859), .B2(n465), .C1(n863), .C2(n485), .A(n759), .ZN(
        n626) );
  AOI22_X1 U627 ( .A1(n870), .A2(a[26]), .B1(a[23]), .B2(n866), .ZN(n759) );
  OAI222_X1 U628 ( .A1(n436), .A2(n308), .B1(n694), .B2(n437), .C1(n438), .C2(
        n343), .ZN(n435) );
  AOI221_X1 U629 ( .B1(a[25]), .B2(n322), .C1(a[28]), .C2(n866), .A(n440), 
        .ZN(n438) );
  AOI222_X1 U630 ( .A1(n310), .A2(n442), .B1(n854), .B2(n443), .C1(n353), .C2(
        n444), .ZN(n437) );
  AOI222_X1 U631 ( .A1(n840), .A2(n445), .B1(n446), .B2(b[3]), .C1(n849), .C2(
        n224), .ZN(n436) );
  OAI222_X1 U632 ( .A1(n415), .A2(n308), .B1(n694), .B2(n416), .C1(n417), .C2(
        n343), .ZN(n414) );
  AOI221_X1 U633 ( .B1(n353), .B2(n192), .C1(n310), .C2(n197), .A(n422), .ZN(
        n415) );
  AOI221_X1 U634 ( .B1(n871), .B2(a[26]), .C1(a[29]), .C2(n866), .A(n418), 
        .ZN(n417) );
  AOI222_X1 U635 ( .A1(n310), .A2(n419), .B1(n854), .B2(n420), .C1(n353), .C2(
        n421), .ZN(n416) );
  OAI222_X1 U636 ( .A1(n376), .A2(n308), .B1(n694), .B2(n377), .C1(n378), .C2(
        n343), .ZN(n375) );
  AOI211_X1 U637 ( .C1(a[28]), .C2(n344), .A(n379), .B(n380), .ZN(n378) );
  AOI221_X1 U638 ( .B1(n310), .B2(n274), .C1(n353), .C2(n275), .A(n386), .ZN(
        n376) );
  AOI222_X1 U639 ( .A1(n310), .A2(n383), .B1(n847), .B2(n384), .C1(n353), .C2(
        n385), .ZN(n377) );
  OAI222_X1 U640 ( .A1(n340), .A2(n308), .B1(n694), .B2(n341), .C1(n342), .C2(
        n343), .ZN(n339) );
  AOI211_X1 U641 ( .C1(n344), .C2(a[29]), .A(n345), .B(n346), .ZN(n342) );
  AOI221_X1 U642 ( .B1(n310), .B2(n256), .C1(n353), .C2(n257), .A(n355), .ZN(
        n340) );
  AOI222_X1 U643 ( .A1(n310), .A2(n350), .B1(n849), .B2(n352), .C1(n353), .C2(
        n354), .ZN(n341) );
  OAI221_X1 U644 ( .B1(n860), .B2(n271), .C1(n325), .C2(n290), .A(n819), .ZN(
        n311) );
  AOI22_X1 U645 ( .A1(a[7]), .A2(n322), .B1(a[4]), .B2(n868), .ZN(n819) );
  AOI21_X1 U646 ( .B1(n834), .B2(a[31]), .A(n380), .ZN(n560) );
  OAI221_X1 U647 ( .B1(n857), .B2(n485), .C1(n864), .C2(n465), .A(n486), .ZN(
        n384) );
  AOI22_X1 U648 ( .A1(a[23]), .A2(n869), .B1(a[26]), .B2(n868), .ZN(n486) );
  OAI221_X1 U649 ( .B1(n857), .B2(n465), .C1(n864), .C2(n441), .A(n466), .ZN(
        n352) );
  AOI22_X1 U650 ( .A1(a[24]), .A2(n869), .B1(a[27]), .B2(n867), .ZN(n466) );
  OAI221_X1 U651 ( .B1(n857), .B2(n248), .C1(n864), .C2(n271), .A(n608), .ZN(
        n291) );
  AOI22_X1 U652 ( .A1(a[8]), .A2(n869), .B1(a[5]), .B2(n868), .ZN(n608) );
  OAI221_X1 U653 ( .B1(n859), .B2(n698), .C1(n862), .C2(n612), .A(n777), .ZN(
        n405) );
  AOI22_X1 U654 ( .A1(a[13]), .A2(n871), .B1(a[10]), .B2(n867), .ZN(n777) );
  OAI221_X1 U655 ( .B1(n859), .B2(n678), .C1(n863), .C2(n698), .A(n762), .ZN(
        n331) );
  AOI22_X1 U656 ( .A1(a[14]), .A2(n871), .B1(a[11]), .B2(n866), .ZN(n762) );
  OAI221_X1 U657 ( .B1(n857), .B2(n522), .C1(n864), .C2(n504), .A(n523), .ZN(
        n443) );
  AOI22_X1 U658 ( .A1(a[21]), .A2(n869), .B1(a[24]), .B2(n867), .ZN(n523) );
  OAI221_X1 U659 ( .B1(n857), .B2(n504), .C1(n864), .C2(n485), .A(n505), .ZN(
        n420) );
  AOI22_X1 U660 ( .A1(a[22]), .A2(n869), .B1(a[25]), .B2(n868), .ZN(n505) );
  OAI221_X1 U661 ( .B1(n858), .B2(n401), .C1(n863), .C2(n328), .A(n738), .ZN(
        n666) );
  AOI22_X1 U662 ( .A1(a[1]), .A2(n871), .B1(a[4]), .B2(n866), .ZN(n738) );
  OAI221_X1 U663 ( .B1(n860), .B2(n641), .C1(n864), .C2(n654), .A(n781), .ZN(
        n402) );
  AOI22_X1 U664 ( .A1(a[17]), .A2(n322), .B1(a[14]), .B2(n867), .ZN(n781) );
  OAI221_X1 U665 ( .B1(n185), .B2(n861), .C1(n325), .C2(n223), .A(n327), .ZN(
        n242) );
  AOI22_X1 U666 ( .A1(a[10]), .A2(n869), .B1(a[7]), .B2(n866), .ZN(n327) );
  OAI221_X1 U667 ( .B1(n185), .B2(n861), .C1(n863), .C2(n613), .A(n763), .ZN(
        n542) );
  AOI22_X1 U668 ( .A1(a[8]), .A2(n871), .B1(a[11]), .B2(n867), .ZN(n763) );
  OAI221_X1 U669 ( .B1(n857), .B2(n223), .C1(n864), .C2(n248), .A(n400), .ZN(
        n265) );
  AOI22_X1 U670 ( .A1(n322), .A2(a[9]), .B1(a[6]), .B2(n868), .ZN(n400) );
  OAI221_X1 U671 ( .B1(n858), .B2(n678), .C1(n325), .C2(n668), .A(n679), .ZN(
        n629) );
  AOI22_X1 U672 ( .A1(a[12]), .A2(n870), .B1(a[15]), .B2(n868), .ZN(n679) );
  AOI22_X1 U673 ( .A1(n737), .A2(n451), .B1(b[2]), .B2(n346), .ZN(n457) );
  AOI221_X1 U674 ( .B1(a[5]), .B2(n322), .C1(a[2]), .C2(n868), .A(n399), .ZN(
        n398) );
  OAI22_X1 U675 ( .A1(n862), .A2(n328), .B1(n861), .B2(n304), .ZN(n399) );
  AOI221_X1 U676 ( .B1(a[6]), .B2(n322), .C1(a[3]), .C2(n867), .A(n324), .ZN(
        n320) );
  OAI22_X1 U677 ( .A1(n862), .A2(n304), .B1(n860), .B2(n290), .ZN(n324) );
  AOI22_X1 U678 ( .A1(n868), .A2(a[1]), .B1(n865), .B2(a[0]), .ZN(n572) );
  OAI221_X1 U679 ( .B1(n349), .B2(n861), .C1(n325), .C2(n382), .A(n814), .ZN(
        n736) );
  AOI22_X1 U680 ( .A1(n870), .A2(a[31]), .B1(a[28]), .B2(n868), .ZN(n814) );
  AOI22_X1 U681 ( .A1(n231), .A2(b[2]), .B1(n737), .B2(n228), .ZN(n446) );
  INV_X1 U682 ( .A(n694), .ZN(n308) );
  AOI21_X1 U683 ( .B1(n865), .B2(a[31]), .A(n380), .ZN(n556) );
  OAI221_X1 U684 ( .B1(n862), .B2(n609), .C1(n872), .C2(n328), .A(n820), .ZN(
        n818) );
  AOI21_X1 U685 ( .B1(a[2]), .B2(n344), .A(n661), .ZN(n820) );
  INV_X1 U686 ( .A(a[27]), .ZN(n381) );
  INV_X1 U687 ( .A(a[24]), .ZN(n485) );
  AOI22_X1 U688 ( .A1(n868), .A2(a[29]), .B1(n865), .B2(a[30]), .ZN(n713) );
  INV_X1 U689 ( .A(b[3]), .ZN(n624) );
  INV_X1 U690 ( .A(a[31]), .ZN(n712) );
  XNOR2_X1 U691 ( .A(n831), .B(a[31]), .ZN(n364) );
  INV_X1 U692 ( .A(a[9]), .ZN(n185) );
  INV_X1 U693 ( .A(a[4]), .ZN(n304) );
  INV_X1 U694 ( .A(a[3]), .ZN(n328) );
  INV_X1 U695 ( .A(a[5]), .ZN(n290) );
  INV_X1 U696 ( .A(a[6]), .ZN(n271) );
  INV_X1 U697 ( .A(a[7]), .ZN(n248) );
  INV_X1 U698 ( .A(a[10]), .ZN(n613) );
  INV_X1 U699 ( .A(a[11]), .ZN(n612) );
  INV_X1 U700 ( .A(a[20]), .ZN(n558) );
  INV_X1 U701 ( .A(a[16]), .ZN(n641) );
  INV_X1 U702 ( .A(a[17]), .ZN(n627) );
  INV_X1 U703 ( .A(a[18]), .ZN(n594) );
  INV_X1 U704 ( .A(a[19]), .ZN(n578) );
  INV_X1 U705 ( .A(a[15]), .ZN(n654) );
  INV_X1 U706 ( .A(a[13]), .ZN(n678) );
  INV_X1 U707 ( .A(a[14]), .ZN(n668) );
  NOR2_X1 U708 ( .A1(n711), .A2(n823), .ZN(n322) );
  INV_X1 U709 ( .A(b[0]), .ZN(n823) );
  INV_X1 U710 ( .A(a[21]), .ZN(n538) );
  NAND2_X1 U711 ( .A1(n310), .A2(a[31]), .ZN(n561) );
  INV_X1 U712 ( .A(a[28]), .ZN(n348) );
  INV_X1 U718 ( .A(a[2]), .ZN(n401) );
  INV_X1 U719 ( .A(a[22]), .ZN(n522) );
  INV_X1 U720 ( .A(a[8]), .ZN(n223) );
  INV_X1 U721 ( .A(a[12]), .ZN(n698) );
  INV_X1 U722 ( .A(b[2]), .ZN(n737) );
  NOR2_X1 U723 ( .A1(n737), .A2(b[3]), .ZN(n351) );
  NOR2_X1 U724 ( .A1(b[3]), .A2(b[2]), .ZN(n439) );
  INV_X1 U725 ( .A(a[30]), .ZN(n349) );
  INV_X1 U726 ( .A(a[29]), .ZN(n382) );
  INV_X1 U727 ( .A(a[26]), .ZN(n441) );
  INV_X1 U728 ( .A(b[1]), .ZN(n711) );
  INV_X1 U729 ( .A(a[25]), .ZN(n465) );
  INV_X1 U730 ( .A(a[23]), .ZN(n504) );
  INV_X1 U731 ( .A(a[1]), .ZN(n609) );
  NAND2_X1 U732 ( .A1(b[0]), .A2(n711), .ZN(n325) );
  INV_X1 U733 ( .A(a[0]), .ZN(n774) );
  OR2_X1 U734 ( .A1(b[0]), .A2(b[1]), .ZN(n834) );
  INV_X1 U735 ( .A(b[6]), .ZN(n269) );
  INV_X1 U736 ( .A(b[7]), .ZN(n246) );
  INV_X1 U737 ( .A(b[22]), .ZN(n552) );
  INV_X1 U738 ( .A(b[31]), .ZN(n831) );
  INV_X1 U739 ( .A(n439), .ZN(n835) );
  INV_X1 U740 ( .A(n439), .ZN(n836) );
  INV_X1 U741 ( .A(n835), .ZN(n837) );
  INV_X1 U742 ( .A(n835), .ZN(n838) );
  INV_X1 U743 ( .A(n835), .ZN(n839) );
  INV_X1 U744 ( .A(n836), .ZN(n840) );
  INV_X1 U745 ( .A(n836), .ZN(n841) );
  INV_X1 U746 ( .A(n836), .ZN(n842) );
  INV_X1 U747 ( .A(n836), .ZN(n843) );
  INV_X1 U748 ( .A(n836), .ZN(n844) );
  INV_X1 U749 ( .A(n351), .ZN(n845) );
  INV_X1 U750 ( .A(n351), .ZN(n846) );
  INV_X1 U751 ( .A(n845), .ZN(n847) );
  INV_X1 U752 ( .A(n845), .ZN(n848) );
  INV_X1 U753 ( .A(n845), .ZN(n849) );
  INV_X1 U754 ( .A(n846), .ZN(n850) );
  INV_X1 U755 ( .A(n846), .ZN(n851) );
  INV_X1 U756 ( .A(n846), .ZN(n852) );
  INV_X1 U757 ( .A(n846), .ZN(n853) );
  INV_X1 U758 ( .A(n846), .ZN(n854) );
  INV_X1 U759 ( .A(n325), .ZN(n865) );
  INV_X1 U760 ( .A(n834), .ZN(n866) );
  INV_X1 U761 ( .A(n834), .ZN(n867) );
  INV_X1 U762 ( .A(n834), .ZN(n868) );
  INV_X1 U763 ( .A(n322), .ZN(n872) );
  INV_X1 U764 ( .A(n189), .ZN(n889) );
  INV_X1 U765 ( .A(n188), .ZN(n892) );
  INV_X1 U766 ( .A(n187), .ZN(n897) );
  INV_X1 U767 ( .A(n187), .ZN(n898) );
  INV_X1 U768 ( .A(n187), .ZN(n899) );
endmodule


module PSWreg ( rst, clk, unaligned, ovf, status );
  output [31:0] status;
  input rst, clk, unaligned, ovf;
  wire   N3, N4, n4;
  assign status[31] = 1'b0;
  assign status[30] = 1'b0;
  assign status[29] = 1'b0;
  assign status[28] = 1'b0;
  assign status[27] = 1'b0;
  assign status[26] = 1'b0;
  assign status[25] = 1'b0;
  assign status[24] = 1'b0;
  assign status[23] = 1'b0;
  assign status[22] = 1'b0;
  assign status[21] = 1'b0;
  assign status[20] = 1'b0;
  assign status[19] = 1'b0;
  assign status[18] = 1'b0;
  assign status[17] = 1'b0;
  assign status[16] = 1'b0;
  assign status[15] = 1'b0;
  assign status[14] = 1'b0;
  assign status[13] = 1'b0;
  assign status[12] = 1'b0;
  assign status[11] = 1'b0;
  assign status[10] = 1'b0;
  assign status[9] = 1'b0;
  assign status[8] = 1'b0;
  assign status[7] = 1'b0;
  assign status[6] = 1'b0;
  assign status[5] = 1'b0;
  assign status[4] = 1'b0;
  assign status[3] = 1'b0;
  assign status[2] = 1'b0;

  DFF_X1 \status_reg[1]  ( .D(N4), .CK(clk), .Q(status[1]) );
  DFF_X1 \status_reg[0]  ( .D(N3), .CK(clk), .Q(status[0]) );
  AND2_X1 U33 ( .A1(unaligned), .A2(n4), .ZN(N3) );
  INV_X1 U34 ( .A(rst), .ZN(n4) );
  AND2_X1 U35 ( .A1(ovf), .A2(n4), .ZN(N4) );
endmodule


module branch_circ ( branch_type, zero, branch_taken );
  input branch_type, zero;
  output branch_taken;


  XOR2_X1 U1 ( .A(zero), .B(branch_type), .Z(branch_taken) );
endmodule


module forward ( rt_addr_IDEX, rs_addr_IDEX, rd_addr_EXMEM, rd_addr_MEMWB, 
        regwrite_EXMEM, regwrite_MEMWB, forwardA, forwardB );
  input [4:0] rt_addr_IDEX;
  input [4:0] rs_addr_IDEX;
  input [4:0] rd_addr_EXMEM;
  input [4:0] rd_addr_MEMWB;
  output [1:0] forwardA;
  output [1:0] forwardB;
  input regwrite_EXMEM, regwrite_MEMWB;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39;

  XOR2_X1 U35 ( .A(rt_addr_IDEX[3]), .B(rd_addr_EXMEM[3]), .Z(n14) );
  XOR2_X1 U36 ( .A(rt_addr_IDEX[2]), .B(rd_addr_EXMEM[2]), .Z(n13) );
  XOR2_X1 U37 ( .A(rt_addr_IDEX[4]), .B(rd_addr_EXMEM[4]), .Z(n12) );
  XOR2_X1 U38 ( .A(rs_addr_IDEX[3]), .B(rd_addr_EXMEM[3]), .Z(n31) );
  XOR2_X1 U39 ( .A(rs_addr_IDEX[2]), .B(rd_addr_EXMEM[2]), .Z(n30) );
  XOR2_X1 U40 ( .A(rs_addr_IDEX[4]), .B(rd_addr_EXMEM[4]), .Z(n29) );
  NOR4_X1 U2 ( .A1(n5), .A2(n6), .A3(forwardB[1]), .A4(n7), .ZN(forwardB[0])
         );
  NAND2_X1 U3 ( .A1(n15), .A2(regwrite_MEMWB), .ZN(n6) );
  NAND4_X1 U4 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n5) );
  XNOR2_X1 U5 ( .A(rd_addr_MEMWB[4]), .B(rt_addr_IDEX[4]), .ZN(n15) );
  NOR4_X1 U6 ( .A1(n20), .A2(n21), .A3(forwardA[1]), .A4(n7), .ZN(forwardA[0])
         );
  NAND2_X1 U7 ( .A1(n35), .A2(regwrite_MEMWB), .ZN(n21) );
  NAND4_X1 U8 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n20) );
  XNOR2_X1 U9 ( .A(rd_addr_MEMWB[4]), .B(rs_addr_IDEX[4]), .ZN(n35) );
  XNOR2_X1 U10 ( .A(rd_addr_MEMWB[2]), .B(rt_addr_IDEX[2]), .ZN(n19) );
  XNOR2_X1 U11 ( .A(rd_addr_MEMWB[2]), .B(rs_addr_IDEX[2]), .ZN(n39) );
  XNOR2_X1 U12 ( .A(rd_addr_MEMWB[1]), .B(rt_addr_IDEX[1]), .ZN(n18) );
  XNOR2_X1 U13 ( .A(rd_addr_MEMWB[0]), .B(rt_addr_IDEX[0]), .ZN(n17) );
  XNOR2_X1 U14 ( .A(rd_addr_MEMWB[1]), .B(rs_addr_IDEX[1]), .ZN(n38) );
  XNOR2_X1 U15 ( .A(rd_addr_MEMWB[0]), .B(rs_addr_IDEX[0]), .ZN(n37) );
  XNOR2_X1 U16 ( .A(rd_addr_MEMWB[3]), .B(rt_addr_IDEX[3]), .ZN(n16) );
  XNOR2_X1 U17 ( .A(rd_addr_MEMWB[3]), .B(rs_addr_IDEX[3]), .ZN(n36) );
  NOR2_X1 U18 ( .A1(rd_addr_MEMWB[1]), .A2(rd_addr_MEMWB[0]), .ZN(n25) );
  AND4_X1 U19 ( .A1(n22), .A2(n23), .A3(n24), .A4(n25), .ZN(n7) );
  INV_X1 U20 ( .A(rd_addr_MEMWB[3]), .ZN(n22) );
  INV_X1 U21 ( .A(rd_addr_MEMWB[4]), .ZN(n23) );
  INV_X1 U22 ( .A(rd_addr_MEMWB[2]), .ZN(n24) );
  INV_X1 U23 ( .A(n32), .ZN(n9) );
  OAI21_X1 U24 ( .B1(n33), .B2(n34), .A(regwrite_EXMEM), .ZN(n32) );
  OR2_X1 U25 ( .A1(rd_addr_EXMEM[0]), .A2(rd_addr_EXMEM[1]), .ZN(n34) );
  OR3_X1 U26 ( .A1(rd_addr_EXMEM[3]), .A2(rd_addr_EXMEM[4]), .A3(
        rd_addr_EXMEM[2]), .ZN(n33) );
  AND4_X1 U27 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(forwardB[1]) );
  XNOR2_X1 U28 ( .A(rd_addr_EXMEM[0]), .B(rt_addr_IDEX[0]), .ZN(n8) );
  XNOR2_X1 U29 ( .A(rd_addr_EXMEM[1]), .B(rt_addr_IDEX[1]), .ZN(n10) );
  NOR3_X1 U30 ( .A1(n12), .A2(n13), .A3(n14), .ZN(n11) );
  AND4_X1 U31 ( .A1(n26), .A2(n9), .A3(n27), .A4(n28), .ZN(forwardA[1]) );
  XNOR2_X1 U32 ( .A(rd_addr_EXMEM[0]), .B(rs_addr_IDEX[0]), .ZN(n26) );
  XNOR2_X1 U33 ( .A(rd_addr_EXMEM[1]), .B(rs_addr_IDEX[1]), .ZN(n27) );
  NOR3_X1 U34 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n28) );
endmodule


module concat16 ( string16, string32 );
  input [15:0] string16;
  output [31:0] string32;
  wire   \string16[15] , \string16[14] , \string16[13] , \string16[12] ,
         \string16[11] , \string16[10] , \string16[9] , \string16[8] ,
         \string16[7] , \string16[6] , \string16[5] , \string16[4] ,
         \string16[3] , \string16[2] , \string16[1] , \string16[0] ;
  assign string32[15] = 1'b0;
  assign string32[14] = 1'b0;
  assign string32[13] = 1'b0;
  assign string32[12] = 1'b0;
  assign string32[11] = 1'b0;
  assign string32[10] = 1'b0;
  assign string32[9] = 1'b0;
  assign string32[8] = 1'b0;
  assign string32[7] = 1'b0;
  assign string32[6] = 1'b0;
  assign string32[5] = 1'b0;
  assign string32[4] = 1'b0;
  assign string32[3] = 1'b0;
  assign string32[2] = 1'b0;
  assign string32[1] = 1'b0;
  assign string32[0] = 1'b0;
  assign string32[31] = \string16[15] ;
  assign \string16[15]  = string16[15];
  assign string32[30] = \string16[14] ;
  assign \string16[14]  = string16[14];
  assign string32[29] = \string16[13] ;
  assign \string16[13]  = string16[13];
  assign string32[28] = \string16[12] ;
  assign \string16[12]  = string16[12];
  assign string32[27] = \string16[11] ;
  assign \string16[11]  = string16[11];
  assign string32[26] = \string16[10] ;
  assign \string16[10]  = string16[10];
  assign string32[25] = \string16[9] ;
  assign \string16[9]  = string16[9];
  assign string32[24] = \string16[8] ;
  assign \string16[8]  = string16[8];
  assign string32[23] = \string16[7] ;
  assign \string16[7]  = string16[7];
  assign string32[22] = \string16[6] ;
  assign \string16[6]  = string16[6];
  assign string32[21] = \string16[5] ;
  assign \string16[5]  = string16[5];
  assign string32[20] = \string16[4] ;
  assign \string16[4]  = string16[4];
  assign string32[19] = \string16[3] ;
  assign \string16[3]  = string16[3];
  assign string32[18] = \string16[2] ;
  assign \string16[2]  = string16[2];
  assign string32[17] = \string16[1] ;
  assign \string16[1]  = string16[1];
  assign string32[16] = \string16[0] ;
  assign \string16[0]  = string16[0];

endmodule


module reg_file ( read_address_1, read_address_2, write_address, write_data, 
        reg_write, rst, data_reg_1, data_reg_2 );
  input [4:0] read_address_1;
  input [4:0] read_address_2;
  input [4:0] write_address;
  input [31:0] write_data;
  output [31:0] data_reg_1;
  output [31:0] data_reg_2;
  input reg_write, rst;
  wire   \bank_register[1][31] , \bank_register[1][30] ,
         \bank_register[1][29] , \bank_register[1][28] ,
         \bank_register[1][27] , \bank_register[1][26] ,
         \bank_register[1][25] , \bank_register[1][24] ,
         \bank_register[1][23] , \bank_register[1][22] ,
         \bank_register[1][21] , \bank_register[1][20] ,
         \bank_register[1][19] , \bank_register[1][18] ,
         \bank_register[1][17] , \bank_register[1][16] ,
         \bank_register[1][15] , \bank_register[1][14] ,
         \bank_register[1][13] , \bank_register[1][12] ,
         \bank_register[1][11] , \bank_register[1][10] , \bank_register[1][9] ,
         \bank_register[1][8] , \bank_register[1][7] , \bank_register[1][6] ,
         \bank_register[1][5] , \bank_register[1][4] , \bank_register[1][3] ,
         \bank_register[1][2] , \bank_register[1][1] , \bank_register[1][0] ,
         \bank_register[2][31] , \bank_register[2][30] ,
         \bank_register[2][29] , \bank_register[2][28] ,
         \bank_register[2][27] , \bank_register[2][26] ,
         \bank_register[2][25] , \bank_register[2][24] ,
         \bank_register[2][23] , \bank_register[2][22] ,
         \bank_register[2][21] , \bank_register[2][20] ,
         \bank_register[2][19] , \bank_register[2][18] ,
         \bank_register[2][17] , \bank_register[2][16] ,
         \bank_register[2][15] , \bank_register[2][14] ,
         \bank_register[2][13] , \bank_register[2][12] ,
         \bank_register[2][11] , \bank_register[2][10] , \bank_register[2][9] ,
         \bank_register[2][8] , \bank_register[2][7] , \bank_register[2][6] ,
         \bank_register[2][5] , \bank_register[2][4] , \bank_register[2][3] ,
         \bank_register[2][2] , \bank_register[2][1] , \bank_register[2][0] ,
         \bank_register[3][31] , \bank_register[3][30] ,
         \bank_register[3][29] , \bank_register[3][28] ,
         \bank_register[3][27] , \bank_register[3][26] ,
         \bank_register[3][25] , \bank_register[3][24] ,
         \bank_register[3][23] , \bank_register[3][22] ,
         \bank_register[3][21] , \bank_register[3][20] ,
         \bank_register[3][19] , \bank_register[3][18] ,
         \bank_register[3][17] , \bank_register[3][16] ,
         \bank_register[3][15] , \bank_register[3][14] ,
         \bank_register[3][13] , \bank_register[3][12] ,
         \bank_register[3][11] , \bank_register[3][10] , \bank_register[3][9] ,
         \bank_register[3][8] , \bank_register[3][7] , \bank_register[3][6] ,
         \bank_register[3][5] , \bank_register[3][4] , \bank_register[3][3] ,
         \bank_register[3][2] , \bank_register[3][1] , \bank_register[3][0] ,
         \bank_register[4][31] , \bank_register[4][30] ,
         \bank_register[4][29] , \bank_register[4][28] ,
         \bank_register[4][27] , \bank_register[4][26] ,
         \bank_register[4][25] , \bank_register[4][24] ,
         \bank_register[4][23] , \bank_register[4][22] ,
         \bank_register[4][21] , \bank_register[4][20] ,
         \bank_register[4][19] , \bank_register[4][18] ,
         \bank_register[4][17] , \bank_register[4][16] ,
         \bank_register[4][15] , \bank_register[4][14] ,
         \bank_register[4][13] , \bank_register[4][12] ,
         \bank_register[4][11] , \bank_register[4][10] , \bank_register[4][9] ,
         \bank_register[4][8] , \bank_register[4][7] , \bank_register[4][6] ,
         \bank_register[4][5] , \bank_register[4][4] , \bank_register[4][3] ,
         \bank_register[4][2] , \bank_register[4][1] , \bank_register[4][0] ,
         \bank_register[5][31] , \bank_register[5][30] ,
         \bank_register[5][29] , \bank_register[5][28] ,
         \bank_register[5][27] , \bank_register[5][26] ,
         \bank_register[5][25] , \bank_register[5][24] ,
         \bank_register[5][23] , \bank_register[5][22] ,
         \bank_register[5][21] , \bank_register[5][20] ,
         \bank_register[5][19] , \bank_register[5][18] ,
         \bank_register[5][17] , \bank_register[5][16] ,
         \bank_register[5][15] , \bank_register[5][14] ,
         \bank_register[5][13] , \bank_register[5][12] ,
         \bank_register[5][11] , \bank_register[5][10] , \bank_register[5][9] ,
         \bank_register[5][8] , \bank_register[5][7] , \bank_register[5][6] ,
         \bank_register[5][5] , \bank_register[5][4] , \bank_register[5][3] ,
         \bank_register[5][2] , \bank_register[5][1] , \bank_register[5][0] ,
         \bank_register[6][31] , \bank_register[6][30] ,
         \bank_register[6][29] , \bank_register[6][28] ,
         \bank_register[6][27] , \bank_register[6][26] ,
         \bank_register[6][25] , \bank_register[6][24] ,
         \bank_register[6][23] , \bank_register[6][22] ,
         \bank_register[6][21] , \bank_register[6][20] ,
         \bank_register[6][19] , \bank_register[6][18] ,
         \bank_register[6][17] , \bank_register[6][16] ,
         \bank_register[6][15] , \bank_register[6][14] ,
         \bank_register[6][13] , \bank_register[6][12] ,
         \bank_register[6][11] , \bank_register[6][10] , \bank_register[6][9] ,
         \bank_register[6][8] , \bank_register[6][7] , \bank_register[6][6] ,
         \bank_register[6][5] , \bank_register[6][4] , \bank_register[6][3] ,
         \bank_register[6][2] , \bank_register[6][1] , \bank_register[6][0] ,
         \bank_register[7][31] , \bank_register[7][30] ,
         \bank_register[7][29] , \bank_register[7][28] ,
         \bank_register[7][27] , \bank_register[7][26] ,
         \bank_register[7][25] , \bank_register[7][24] ,
         \bank_register[7][23] , \bank_register[7][22] ,
         \bank_register[7][21] , \bank_register[7][20] ,
         \bank_register[7][19] , \bank_register[7][18] ,
         \bank_register[7][17] , \bank_register[7][16] ,
         \bank_register[7][15] , \bank_register[7][14] ,
         \bank_register[7][13] , \bank_register[7][12] ,
         \bank_register[7][11] , \bank_register[7][10] , \bank_register[7][9] ,
         \bank_register[7][8] , \bank_register[7][7] , \bank_register[7][6] ,
         \bank_register[7][5] , \bank_register[7][4] , \bank_register[7][3] ,
         \bank_register[7][2] , \bank_register[7][1] , \bank_register[7][0] ,
         \bank_register[8][31] , \bank_register[8][30] ,
         \bank_register[8][29] , \bank_register[8][28] ,
         \bank_register[8][27] , \bank_register[8][26] ,
         \bank_register[8][25] , \bank_register[8][24] ,
         \bank_register[8][23] , \bank_register[8][22] ,
         \bank_register[8][21] , \bank_register[8][20] ,
         \bank_register[8][19] , \bank_register[8][18] ,
         \bank_register[8][17] , \bank_register[8][16] ,
         \bank_register[8][15] , \bank_register[8][14] ,
         \bank_register[8][13] , \bank_register[8][12] ,
         \bank_register[8][11] , \bank_register[8][10] , \bank_register[8][9] ,
         \bank_register[8][8] , \bank_register[8][7] , \bank_register[8][6] ,
         \bank_register[8][5] , \bank_register[8][4] , \bank_register[8][3] ,
         \bank_register[8][2] , \bank_register[8][1] , \bank_register[8][0] ,
         \bank_register[9][31] , \bank_register[9][30] ,
         \bank_register[9][29] , \bank_register[9][28] ,
         \bank_register[9][27] , \bank_register[9][26] ,
         \bank_register[9][25] , \bank_register[9][24] ,
         \bank_register[9][23] , \bank_register[9][22] ,
         \bank_register[9][21] , \bank_register[9][20] ,
         \bank_register[9][19] , \bank_register[9][18] ,
         \bank_register[9][17] , \bank_register[9][16] ,
         \bank_register[9][15] , \bank_register[9][14] ,
         \bank_register[9][13] , \bank_register[9][12] ,
         \bank_register[9][11] , \bank_register[9][10] , \bank_register[9][9] ,
         \bank_register[9][8] , \bank_register[9][7] , \bank_register[9][6] ,
         \bank_register[9][5] , \bank_register[9][4] , \bank_register[9][3] ,
         \bank_register[9][2] , \bank_register[9][1] , \bank_register[9][0] ,
         \bank_register[10][31] , \bank_register[10][30] ,
         \bank_register[10][29] , \bank_register[10][28] ,
         \bank_register[10][27] , \bank_register[10][26] ,
         \bank_register[10][25] , \bank_register[10][24] ,
         \bank_register[10][23] , \bank_register[10][22] ,
         \bank_register[10][21] , \bank_register[10][20] ,
         \bank_register[10][19] , \bank_register[10][18] ,
         \bank_register[10][17] , \bank_register[10][16] ,
         \bank_register[10][15] , \bank_register[10][14] ,
         \bank_register[10][13] , \bank_register[10][12] ,
         \bank_register[10][11] , \bank_register[10][10] ,
         \bank_register[10][9] , \bank_register[10][8] ,
         \bank_register[10][7] , \bank_register[10][6] ,
         \bank_register[10][5] , \bank_register[10][4] ,
         \bank_register[10][3] , \bank_register[10][2] ,
         \bank_register[10][1] , \bank_register[10][0] ,
         \bank_register[11][31] , \bank_register[11][30] ,
         \bank_register[11][29] , \bank_register[11][28] ,
         \bank_register[11][27] , \bank_register[11][26] ,
         \bank_register[11][25] , \bank_register[11][24] ,
         \bank_register[11][23] , \bank_register[11][22] ,
         \bank_register[11][21] , \bank_register[11][20] ,
         \bank_register[11][19] , \bank_register[11][18] ,
         \bank_register[11][17] , \bank_register[11][16] ,
         \bank_register[11][15] , \bank_register[11][14] ,
         \bank_register[11][13] , \bank_register[11][12] ,
         \bank_register[11][11] , \bank_register[11][10] ,
         \bank_register[11][9] , \bank_register[11][8] ,
         \bank_register[11][7] , \bank_register[11][6] ,
         \bank_register[11][5] , \bank_register[11][4] ,
         \bank_register[11][3] , \bank_register[11][2] ,
         \bank_register[11][1] , \bank_register[11][0] ,
         \bank_register[12][31] , \bank_register[12][30] ,
         \bank_register[12][29] , \bank_register[12][28] ,
         \bank_register[12][27] , \bank_register[12][26] ,
         \bank_register[12][25] , \bank_register[12][24] ,
         \bank_register[12][23] , \bank_register[12][22] ,
         \bank_register[12][21] , \bank_register[12][20] ,
         \bank_register[12][19] , \bank_register[12][18] ,
         \bank_register[12][17] , \bank_register[12][16] ,
         \bank_register[12][15] , \bank_register[12][14] ,
         \bank_register[12][13] , \bank_register[12][12] ,
         \bank_register[12][11] , \bank_register[12][10] ,
         \bank_register[12][9] , \bank_register[12][8] ,
         \bank_register[12][7] , \bank_register[12][6] ,
         \bank_register[12][5] , \bank_register[12][4] ,
         \bank_register[12][3] , \bank_register[12][2] ,
         \bank_register[12][1] , \bank_register[12][0] ,
         \bank_register[13][31] , \bank_register[13][30] ,
         \bank_register[13][29] , \bank_register[13][28] ,
         \bank_register[13][27] , \bank_register[13][26] ,
         \bank_register[13][25] , \bank_register[13][24] ,
         \bank_register[13][23] , \bank_register[13][22] ,
         \bank_register[13][21] , \bank_register[13][20] ,
         \bank_register[13][19] , \bank_register[13][18] ,
         \bank_register[13][17] , \bank_register[13][16] ,
         \bank_register[13][15] , \bank_register[13][14] ,
         \bank_register[13][13] , \bank_register[13][12] ,
         \bank_register[13][11] , \bank_register[13][10] ,
         \bank_register[13][9] , \bank_register[13][8] ,
         \bank_register[13][7] , \bank_register[13][6] ,
         \bank_register[13][5] , \bank_register[13][4] ,
         \bank_register[13][3] , \bank_register[13][2] ,
         \bank_register[13][1] , \bank_register[13][0] ,
         \bank_register[14][31] , \bank_register[14][30] ,
         \bank_register[14][29] , \bank_register[14][28] ,
         \bank_register[14][27] , \bank_register[14][26] ,
         \bank_register[14][25] , \bank_register[14][24] ,
         \bank_register[14][23] , \bank_register[14][22] ,
         \bank_register[14][21] , \bank_register[14][20] ,
         \bank_register[14][19] , \bank_register[14][18] ,
         \bank_register[14][17] , \bank_register[14][16] ,
         \bank_register[14][15] , \bank_register[14][14] ,
         \bank_register[14][13] , \bank_register[14][12] ,
         \bank_register[14][11] , \bank_register[14][10] ,
         \bank_register[14][9] , \bank_register[14][8] ,
         \bank_register[14][7] , \bank_register[14][6] ,
         \bank_register[14][5] , \bank_register[14][4] ,
         \bank_register[14][3] , \bank_register[14][2] ,
         \bank_register[14][1] , \bank_register[14][0] ,
         \bank_register[15][31] , \bank_register[15][30] ,
         \bank_register[15][29] , \bank_register[15][28] ,
         \bank_register[15][27] , \bank_register[15][26] ,
         \bank_register[15][25] , \bank_register[15][24] ,
         \bank_register[15][23] , \bank_register[15][22] ,
         \bank_register[15][21] , \bank_register[15][20] ,
         \bank_register[15][19] , \bank_register[15][18] ,
         \bank_register[15][17] , \bank_register[15][16] ,
         \bank_register[15][15] , \bank_register[15][14] ,
         \bank_register[15][13] , \bank_register[15][12] ,
         \bank_register[15][11] , \bank_register[15][10] ,
         \bank_register[15][9] , \bank_register[15][8] ,
         \bank_register[15][7] , \bank_register[15][6] ,
         \bank_register[15][5] , \bank_register[15][4] ,
         \bank_register[15][3] , \bank_register[15][2] ,
         \bank_register[15][1] , \bank_register[15][0] ,
         \bank_register[16][31] , \bank_register[16][30] ,
         \bank_register[16][29] , \bank_register[16][28] ,
         \bank_register[16][27] , \bank_register[16][26] ,
         \bank_register[16][25] , \bank_register[16][24] ,
         \bank_register[16][23] , \bank_register[16][22] ,
         \bank_register[16][21] , \bank_register[16][20] ,
         \bank_register[16][19] , \bank_register[16][18] ,
         \bank_register[16][17] , \bank_register[16][16] ,
         \bank_register[16][15] , \bank_register[16][14] ,
         \bank_register[16][13] , \bank_register[16][12] ,
         \bank_register[16][11] , \bank_register[16][10] ,
         \bank_register[16][9] , \bank_register[16][8] ,
         \bank_register[16][7] , \bank_register[16][6] ,
         \bank_register[16][5] , \bank_register[16][4] ,
         \bank_register[16][3] , \bank_register[16][2] ,
         \bank_register[16][1] , \bank_register[16][0] ,
         \bank_register[17][31] , \bank_register[17][30] ,
         \bank_register[17][29] , \bank_register[17][28] ,
         \bank_register[17][27] , \bank_register[17][26] ,
         \bank_register[17][25] , \bank_register[17][24] ,
         \bank_register[17][23] , \bank_register[17][22] ,
         \bank_register[17][21] , \bank_register[17][20] ,
         \bank_register[17][19] , \bank_register[17][18] ,
         \bank_register[17][17] , \bank_register[17][16] ,
         \bank_register[17][15] , \bank_register[17][14] ,
         \bank_register[17][13] , \bank_register[17][12] ,
         \bank_register[17][11] , \bank_register[17][10] ,
         \bank_register[17][9] , \bank_register[17][8] ,
         \bank_register[17][7] , \bank_register[17][6] ,
         \bank_register[17][5] , \bank_register[17][4] ,
         \bank_register[17][3] , \bank_register[17][2] ,
         \bank_register[17][1] , \bank_register[17][0] ,
         \bank_register[18][31] , \bank_register[18][30] ,
         \bank_register[18][29] , \bank_register[18][28] ,
         \bank_register[18][27] , \bank_register[18][26] ,
         \bank_register[18][25] , \bank_register[18][24] ,
         \bank_register[18][23] , \bank_register[18][22] ,
         \bank_register[18][21] , \bank_register[18][20] ,
         \bank_register[18][19] , \bank_register[18][18] ,
         \bank_register[18][17] , \bank_register[18][16] ,
         \bank_register[18][15] , \bank_register[18][14] ,
         \bank_register[18][13] , \bank_register[18][12] ,
         \bank_register[18][11] , \bank_register[18][10] ,
         \bank_register[18][9] , \bank_register[18][8] ,
         \bank_register[18][7] , \bank_register[18][6] ,
         \bank_register[18][5] , \bank_register[18][4] ,
         \bank_register[18][3] , \bank_register[18][2] ,
         \bank_register[18][1] , \bank_register[18][0] ,
         \bank_register[19][31] , \bank_register[19][30] ,
         \bank_register[19][29] , \bank_register[19][28] ,
         \bank_register[19][27] , \bank_register[19][26] ,
         \bank_register[19][25] , \bank_register[19][24] ,
         \bank_register[19][23] , \bank_register[19][22] ,
         \bank_register[19][21] , \bank_register[19][20] ,
         \bank_register[19][19] , \bank_register[19][18] ,
         \bank_register[19][17] , \bank_register[19][16] ,
         \bank_register[19][15] , \bank_register[19][14] ,
         \bank_register[19][13] , \bank_register[19][12] ,
         \bank_register[19][11] , \bank_register[19][10] ,
         \bank_register[19][9] , \bank_register[19][8] ,
         \bank_register[19][7] , \bank_register[19][6] ,
         \bank_register[19][5] , \bank_register[19][4] ,
         \bank_register[19][3] , \bank_register[19][2] ,
         \bank_register[19][1] , \bank_register[19][0] ,
         \bank_register[20][31] , \bank_register[20][30] ,
         \bank_register[20][29] , \bank_register[20][28] ,
         \bank_register[20][27] , \bank_register[20][26] ,
         \bank_register[20][25] , \bank_register[20][24] ,
         \bank_register[20][23] , \bank_register[20][22] ,
         \bank_register[20][21] , \bank_register[20][20] ,
         \bank_register[20][19] , \bank_register[20][18] ,
         \bank_register[20][17] , \bank_register[20][16] ,
         \bank_register[20][15] , \bank_register[20][14] ,
         \bank_register[20][13] , \bank_register[20][12] ,
         \bank_register[20][11] , \bank_register[20][10] ,
         \bank_register[20][9] , \bank_register[20][8] ,
         \bank_register[20][7] , \bank_register[20][6] ,
         \bank_register[20][5] , \bank_register[20][4] ,
         \bank_register[20][3] , \bank_register[20][2] ,
         \bank_register[20][1] , \bank_register[20][0] ,
         \bank_register[21][31] , \bank_register[21][30] ,
         \bank_register[21][29] , \bank_register[21][28] ,
         \bank_register[21][27] , \bank_register[21][26] ,
         \bank_register[21][25] , \bank_register[21][24] ,
         \bank_register[21][23] , \bank_register[21][22] ,
         \bank_register[21][21] , \bank_register[21][20] ,
         \bank_register[21][19] , \bank_register[21][18] ,
         \bank_register[21][17] , \bank_register[21][16] ,
         \bank_register[21][15] , \bank_register[21][14] ,
         \bank_register[21][13] , \bank_register[21][12] ,
         \bank_register[21][11] , \bank_register[21][10] ,
         \bank_register[21][9] , \bank_register[21][8] ,
         \bank_register[21][7] , \bank_register[21][6] ,
         \bank_register[21][5] , \bank_register[21][4] ,
         \bank_register[21][3] , \bank_register[21][2] ,
         \bank_register[21][1] , \bank_register[21][0] ,
         \bank_register[22][31] , \bank_register[22][30] ,
         \bank_register[22][29] , \bank_register[22][28] ,
         \bank_register[22][27] , \bank_register[22][26] ,
         \bank_register[22][25] , \bank_register[22][24] ,
         \bank_register[22][23] , \bank_register[22][22] ,
         \bank_register[22][21] , \bank_register[22][20] ,
         \bank_register[22][19] , \bank_register[22][18] ,
         \bank_register[22][17] , \bank_register[22][16] ,
         \bank_register[22][15] , \bank_register[22][14] ,
         \bank_register[22][13] , \bank_register[22][12] ,
         \bank_register[22][11] , \bank_register[22][10] ,
         \bank_register[22][9] , \bank_register[22][8] ,
         \bank_register[22][7] , \bank_register[22][6] ,
         \bank_register[22][5] , \bank_register[22][4] ,
         \bank_register[22][3] , \bank_register[22][2] ,
         \bank_register[22][1] , \bank_register[22][0] ,
         \bank_register[23][31] , \bank_register[23][30] ,
         \bank_register[23][29] , \bank_register[23][28] ,
         \bank_register[23][27] , \bank_register[23][26] ,
         \bank_register[23][25] , \bank_register[23][24] ,
         \bank_register[23][23] , \bank_register[23][22] ,
         \bank_register[23][21] , \bank_register[23][20] ,
         \bank_register[23][19] , \bank_register[23][18] ,
         \bank_register[23][17] , \bank_register[23][16] ,
         \bank_register[23][15] , \bank_register[23][14] ,
         \bank_register[23][13] , \bank_register[23][12] ,
         \bank_register[23][11] , \bank_register[23][10] ,
         \bank_register[23][9] , \bank_register[23][8] ,
         \bank_register[23][7] , \bank_register[23][6] ,
         \bank_register[23][5] , \bank_register[23][4] ,
         \bank_register[23][3] , \bank_register[23][2] ,
         \bank_register[23][1] , \bank_register[23][0] ,
         \bank_register[24][31] , \bank_register[24][30] ,
         \bank_register[24][29] , \bank_register[24][28] ,
         \bank_register[24][27] , \bank_register[24][26] ,
         \bank_register[24][25] , \bank_register[24][24] ,
         \bank_register[24][23] , \bank_register[24][22] ,
         \bank_register[24][21] , \bank_register[24][20] ,
         \bank_register[24][19] , \bank_register[24][18] ,
         \bank_register[24][17] , \bank_register[24][16] ,
         \bank_register[24][15] , \bank_register[24][14] ,
         \bank_register[24][13] , \bank_register[24][12] ,
         \bank_register[24][11] , \bank_register[24][10] ,
         \bank_register[24][9] , \bank_register[24][8] ,
         \bank_register[24][7] , \bank_register[24][6] ,
         \bank_register[24][5] , \bank_register[24][4] ,
         \bank_register[24][3] , \bank_register[24][2] ,
         \bank_register[24][1] , \bank_register[24][0] ,
         \bank_register[25][31] , \bank_register[25][30] ,
         \bank_register[25][29] , \bank_register[25][28] ,
         \bank_register[25][27] , \bank_register[25][26] ,
         \bank_register[25][25] , \bank_register[25][24] ,
         \bank_register[25][23] , \bank_register[25][22] ,
         \bank_register[25][21] , \bank_register[25][20] ,
         \bank_register[25][19] , \bank_register[25][18] ,
         \bank_register[25][17] , \bank_register[25][16] ,
         \bank_register[25][15] , \bank_register[25][14] ,
         \bank_register[25][13] , \bank_register[25][12] ,
         \bank_register[25][11] , \bank_register[25][10] ,
         \bank_register[25][9] , \bank_register[25][8] ,
         \bank_register[25][7] , \bank_register[25][6] ,
         \bank_register[25][5] , \bank_register[25][4] ,
         \bank_register[25][3] , \bank_register[25][2] ,
         \bank_register[25][1] , \bank_register[25][0] ,
         \bank_register[26][31] , \bank_register[26][30] ,
         \bank_register[26][29] , \bank_register[26][28] ,
         \bank_register[26][27] , \bank_register[26][26] ,
         \bank_register[26][25] , \bank_register[26][24] ,
         \bank_register[26][23] , \bank_register[26][22] ,
         \bank_register[26][21] , \bank_register[26][20] ,
         \bank_register[26][19] , \bank_register[26][18] ,
         \bank_register[26][17] , \bank_register[26][16] ,
         \bank_register[26][15] , \bank_register[26][14] ,
         \bank_register[26][13] , \bank_register[26][12] ,
         \bank_register[26][11] , \bank_register[26][10] ,
         \bank_register[26][9] , \bank_register[26][8] ,
         \bank_register[26][7] , \bank_register[26][6] ,
         \bank_register[26][5] , \bank_register[26][4] ,
         \bank_register[26][3] , \bank_register[26][2] ,
         \bank_register[26][1] , \bank_register[26][0] ,
         \bank_register[27][31] , \bank_register[27][30] ,
         \bank_register[27][29] , \bank_register[27][28] ,
         \bank_register[27][27] , \bank_register[27][26] ,
         \bank_register[27][25] , \bank_register[27][24] ,
         \bank_register[27][23] , \bank_register[27][22] ,
         \bank_register[27][21] , \bank_register[27][20] ,
         \bank_register[27][19] , \bank_register[27][18] ,
         \bank_register[27][17] , \bank_register[27][16] ,
         \bank_register[27][15] , \bank_register[27][14] ,
         \bank_register[27][13] , \bank_register[27][12] ,
         \bank_register[27][11] , \bank_register[27][10] ,
         \bank_register[27][9] , \bank_register[27][8] ,
         \bank_register[27][7] , \bank_register[27][6] ,
         \bank_register[27][5] , \bank_register[27][4] ,
         \bank_register[27][3] , \bank_register[27][2] ,
         \bank_register[27][1] , \bank_register[27][0] ,
         \bank_register[28][31] , \bank_register[28][30] ,
         \bank_register[28][29] , \bank_register[28][28] ,
         \bank_register[28][27] , \bank_register[28][26] ,
         \bank_register[28][25] , \bank_register[28][24] ,
         \bank_register[28][23] , \bank_register[28][22] ,
         \bank_register[28][21] , \bank_register[28][20] ,
         \bank_register[28][19] , \bank_register[28][18] ,
         \bank_register[28][17] , \bank_register[28][16] ,
         \bank_register[28][15] , \bank_register[28][14] ,
         \bank_register[28][13] , \bank_register[28][12] ,
         \bank_register[28][11] , \bank_register[28][10] ,
         \bank_register[28][9] , \bank_register[28][8] ,
         \bank_register[28][7] , \bank_register[28][6] ,
         \bank_register[28][5] , \bank_register[28][4] ,
         \bank_register[28][3] , \bank_register[28][2] ,
         \bank_register[28][1] , \bank_register[28][0] ,
         \bank_register[29][31] , \bank_register[29][30] ,
         \bank_register[29][29] , \bank_register[29][28] ,
         \bank_register[29][27] , \bank_register[29][26] ,
         \bank_register[29][25] , \bank_register[29][24] ,
         \bank_register[29][23] , \bank_register[29][22] ,
         \bank_register[29][21] , \bank_register[29][20] ,
         \bank_register[29][19] , \bank_register[29][18] ,
         \bank_register[29][17] , \bank_register[29][16] ,
         \bank_register[29][15] , \bank_register[29][14] ,
         \bank_register[29][13] , \bank_register[29][12] ,
         \bank_register[29][11] , \bank_register[29][10] ,
         \bank_register[29][9] , \bank_register[29][8] ,
         \bank_register[29][7] , \bank_register[29][6] ,
         \bank_register[29][5] , \bank_register[29][4] ,
         \bank_register[29][3] , \bank_register[29][2] ,
         \bank_register[29][1] , \bank_register[29][0] ,
         \bank_register[30][31] , \bank_register[30][30] ,
         \bank_register[30][29] , \bank_register[30][28] ,
         \bank_register[30][27] , \bank_register[30][26] ,
         \bank_register[30][25] , \bank_register[30][24] ,
         \bank_register[30][23] , \bank_register[30][22] ,
         \bank_register[30][21] , \bank_register[30][20] ,
         \bank_register[30][19] , \bank_register[30][18] ,
         \bank_register[30][17] , \bank_register[30][16] ,
         \bank_register[30][15] , \bank_register[30][14] ,
         \bank_register[30][13] , \bank_register[30][12] ,
         \bank_register[30][11] , \bank_register[30][10] ,
         \bank_register[30][9] , \bank_register[30][8] ,
         \bank_register[30][7] , \bank_register[30][6] ,
         \bank_register[30][5] , \bank_register[30][4] ,
         \bank_register[30][3] , \bank_register[30][2] ,
         \bank_register[30][1] , \bank_register[30][0] ,
         \bank_register[31][31] , \bank_register[31][30] ,
         \bank_register[31][29] , \bank_register[31][28] ,
         \bank_register[31][27] , \bank_register[31][26] ,
         \bank_register[31][25] , \bank_register[31][24] ,
         \bank_register[31][23] , \bank_register[31][22] ,
         \bank_register[31][21] , \bank_register[31][20] ,
         \bank_register[31][19] , \bank_register[31][18] ,
         \bank_register[31][17] , \bank_register[31][16] ,
         \bank_register[31][15] , \bank_register[31][14] ,
         \bank_register[31][13] , \bank_register[31][12] ,
         \bank_register[31][11] , \bank_register[31][10] ,
         \bank_register[31][9] , \bank_register[31][8] ,
         \bank_register[31][7] , \bank_register[31][6] ,
         \bank_register[31][5] , \bank_register[31][4] ,
         \bank_register[31][3] , \bank_register[31][2] ,
         \bank_register[31][1] , \bank_register[31][0] , N4144, n2152, n2155,
         n2158, n2161, n2164, n2167, n2170, n2173, n2176, n2179, n2182, n2185,
         n2188, n2191, n2194, n2197, n2200, n2203, n2206, n2209, n2212, n2215,
         n2218, n2221, n2224, n2227, n2230, n2233, n2236, n2239, n2242, n2245,
         n2249, n2253, n2257, n2261, n2265, n2269, n2273, n2277, n2281, n2285,
         n2289, n2293, n2297, n2301, n2305, n2309, n2313, n2317, n2321, n2325,
         n2329, n2333, n2337, n2341, n2345, n2349, n2353, n2357, n2361, n2365,
         n2369, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2153,
         n2154, n2156, n2157, n2159, n2160, n2162, n2163, n2165, n2166, n2168,
         n2169, n2171, n2172, n2174, n2175, n2177, n2178, n2180, n2181, n2183,
         n2184, n2186, n2187, n2189, n2190, n2192, n2193, n2195, n2196, n2198,
         n2199, n2201, n2202, n2204, n2205, n2207, n2208, n2210, n2211, n2213,
         n2214, n2216, n2217, n2219, n2220, n2222, n2223, n2225, n2226, n2228,
         n2229, n2231, n2232, n2234, n2235, n2237, n2238, n2240, n2241, n2243,
         n2244, n2246, n2247, n2248, n2250, n2251, n2252, n2254, n2255, n2256,
         n2258, n2259, n2260, n2262, n2263, n2264, n2266, n2267, n2268, n2270,
         n2271, n2272, n2274, n2275, n2276, n2278, n2279, n2280, n2282, n2283,
         n2284, n2286, n2287, n2288, n2290, n2291, n2292, n2294, n2295, n2296,
         n2298, n2299, n2300, n2302, n2303, n2304, n2306, n2307, n2308, n2310,
         n2311, n2312, n2314, n2315, n2316, n2318, n2319, n2320, n2322, n2323,
         n2324, n2326, n2327, n2328, n2330, n2331, n2332, n2334, n2335, n2336,
         n2338, n2339, n2340, n2342, n2343, n2344, n2346, n2347, n2348, n2350,
         n2351, n2352, n2354, n2355, n2356, n2358, n2359, n2360, n2362, n2363,
         n2364, n2366, n2367, n2368, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2767, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241;
  assign N4144 = rst;

  DLH_X1 \bank_register_reg[1][31]  ( .G(n3141), .D(n3235), .Q(
        \bank_register[1][31] ) );
  DLH_X1 \bank_register_reg[1][30]  ( .G(n3141), .D(n3232), .Q(
        \bank_register[1][30] ) );
  DLH_X1 \bank_register_reg[1][29]  ( .G(n3139), .D(n3229), .Q(
        \bank_register[1][29] ) );
  DLH_X1 \bank_register_reg[1][28]  ( .G(n3139), .D(n3226), .Q(
        \bank_register[1][28] ) );
  DLH_X1 \bank_register_reg[1][27]  ( .G(n3139), .D(n3223), .Q(
        \bank_register[1][27] ) );
  DLH_X1 \bank_register_reg[1][26]  ( .G(n3139), .D(n3220), .Q(
        \bank_register[1][26] ) );
  DLH_X1 \bank_register_reg[1][25]  ( .G(n3139), .D(n3217), .Q(
        \bank_register[1][25] ) );
  DLH_X1 \bank_register_reg[1][24]  ( .G(n3139), .D(n3214), .Q(
        \bank_register[1][24] ) );
  DLH_X1 \bank_register_reg[1][23]  ( .G(n3139), .D(n3211), .Q(
        \bank_register[1][23] ) );
  DLH_X1 \bank_register_reg[1][22]  ( .G(n3139), .D(n3208), .Q(
        \bank_register[1][22] ) );
  DLH_X1 \bank_register_reg[1][21]  ( .G(n3139), .D(n3205), .Q(
        \bank_register[1][21] ) );
  DLH_X1 \bank_register_reg[1][20]  ( .G(n3139), .D(n3202), .Q(
        \bank_register[1][20] ) );
  DLH_X1 \bank_register_reg[1][19]  ( .G(n3140), .D(n3199), .Q(
        \bank_register[1][19] ) );
  DLH_X1 \bank_register_reg[1][18]  ( .G(n3140), .D(n3196), .Q(
        \bank_register[1][18] ) );
  DLH_X1 \bank_register_reg[1][17]  ( .G(n3141), .D(n3193), .Q(
        \bank_register[1][17] ) );
  DLH_X1 \bank_register_reg[1][16]  ( .G(n3141), .D(n3190), .Q(
        \bank_register[1][16] ) );
  DLH_X1 \bank_register_reg[1][15]  ( .G(n3141), .D(n3187), .Q(
        \bank_register[1][15] ) );
  DLH_X1 \bank_register_reg[1][14]  ( .G(n3141), .D(n3184), .Q(
        \bank_register[1][14] ) );
  DLH_X1 \bank_register_reg[1][13]  ( .G(n3141), .D(n3181), .Q(
        \bank_register[1][13] ) );
  DLH_X1 \bank_register_reg[1][12]  ( .G(n3141), .D(n3178), .Q(
        \bank_register[1][12] ) );
  DLH_X1 \bank_register_reg[1][11]  ( .G(n3141), .D(n3175), .Q(
        \bank_register[1][11] ) );
  DLH_X1 \bank_register_reg[1][10]  ( .G(n3141), .D(n3172), .Q(
        \bank_register[1][10] ) );
  DLH_X1 \bank_register_reg[1][9]  ( .G(n3140), .D(n3169), .Q(
        \bank_register[1][9] ) );
  DLH_X1 \bank_register_reg[1][8]  ( .G(n3140), .D(n3166), .Q(
        \bank_register[1][8] ) );
  DLH_X1 \bank_register_reg[1][7]  ( .G(n3140), .D(n3163), .Q(
        \bank_register[1][7] ) );
  DLH_X1 \bank_register_reg[1][6]  ( .G(n3140), .D(n3160), .Q(
        \bank_register[1][6] ) );
  DLH_X1 \bank_register_reg[1][5]  ( .G(n3140), .D(n3157), .Q(
        \bank_register[1][5] ) );
  DLH_X1 \bank_register_reg[1][4]  ( .G(n3140), .D(n3154), .Q(
        \bank_register[1][4] ) );
  DLH_X1 \bank_register_reg[1][3]  ( .G(n3140), .D(n3151), .Q(
        \bank_register[1][3] ) );
  DLH_X1 \bank_register_reg[1][2]  ( .G(n3140), .D(n3148), .Q(
        \bank_register[1][2] ) );
  DLH_X1 \bank_register_reg[1][1]  ( .G(n3140), .D(n3145), .Q(
        \bank_register[1][1] ) );
  DLH_X1 \bank_register_reg[1][0]  ( .G(n3139), .D(n3142), .Q(
        \bank_register[1][0] ) );
  DLH_X1 \bank_register_reg[2][31]  ( .G(n3138), .D(n3236), .Q(
        \bank_register[2][31] ) );
  DLH_X1 \bank_register_reg[2][30]  ( .G(n3138), .D(n3233), .Q(
        \bank_register[2][30] ) );
  DLH_X1 \bank_register_reg[2][29]  ( .G(n3136), .D(n3230), .Q(
        \bank_register[2][29] ) );
  DLH_X1 \bank_register_reg[2][28]  ( .G(n3136), .D(n3227), .Q(
        \bank_register[2][28] ) );
  DLH_X1 \bank_register_reg[2][27]  ( .G(n3136), .D(n3224), .Q(
        \bank_register[2][27] ) );
  DLH_X1 \bank_register_reg[2][26]  ( .G(n3136), .D(n3221), .Q(
        \bank_register[2][26] ) );
  DLH_X1 \bank_register_reg[2][25]  ( .G(n3136), .D(n3218), .Q(
        \bank_register[2][25] ) );
  DLH_X1 \bank_register_reg[2][24]  ( .G(n3136), .D(n3215), .Q(
        \bank_register[2][24] ) );
  DLH_X1 \bank_register_reg[2][23]  ( .G(n3136), .D(n3212), .Q(
        \bank_register[2][23] ) );
  DLH_X1 \bank_register_reg[2][22]  ( .G(n3136), .D(n3209), .Q(
        \bank_register[2][22] ) );
  DLH_X1 \bank_register_reg[2][21]  ( .G(n3136), .D(n3206), .Q(
        \bank_register[2][21] ) );
  DLH_X1 \bank_register_reg[2][20]  ( .G(n3136), .D(n3203), .Q(
        \bank_register[2][20] ) );
  DLH_X1 \bank_register_reg[2][19]  ( .G(n3137), .D(n3200), .Q(
        \bank_register[2][19] ) );
  DLH_X1 \bank_register_reg[2][18]  ( .G(n3137), .D(n3197), .Q(
        \bank_register[2][18] ) );
  DLH_X1 \bank_register_reg[2][17]  ( .G(n3138), .D(n3194), .Q(
        \bank_register[2][17] ) );
  DLH_X1 \bank_register_reg[2][16]  ( .G(n3138), .D(n3191), .Q(
        \bank_register[2][16] ) );
  DLH_X1 \bank_register_reg[2][15]  ( .G(n3138), .D(n3188), .Q(
        \bank_register[2][15] ) );
  DLH_X1 \bank_register_reg[2][14]  ( .G(n3138), .D(n3185), .Q(
        \bank_register[2][14] ) );
  DLH_X1 \bank_register_reg[2][13]  ( .G(n3138), .D(n3182), .Q(
        \bank_register[2][13] ) );
  DLH_X1 \bank_register_reg[2][12]  ( .G(n3138), .D(n3179), .Q(
        \bank_register[2][12] ) );
  DLH_X1 \bank_register_reg[2][11]  ( .G(n3138), .D(n3176), .Q(
        \bank_register[2][11] ) );
  DLH_X1 \bank_register_reg[2][10]  ( .G(n3138), .D(n3173), .Q(
        \bank_register[2][10] ) );
  DLH_X1 \bank_register_reg[2][9]  ( .G(n3137), .D(n3170), .Q(
        \bank_register[2][9] ) );
  DLH_X1 \bank_register_reg[2][8]  ( .G(n3137), .D(n3167), .Q(
        \bank_register[2][8] ) );
  DLH_X1 \bank_register_reg[2][7]  ( .G(n3137), .D(n3164), .Q(
        \bank_register[2][7] ) );
  DLH_X1 \bank_register_reg[2][6]  ( .G(n3137), .D(n3161), .Q(
        \bank_register[2][6] ) );
  DLH_X1 \bank_register_reg[2][5]  ( .G(n3137), .D(n3158), .Q(
        \bank_register[2][5] ) );
  DLH_X1 \bank_register_reg[2][4]  ( .G(n3137), .D(n3155), .Q(
        \bank_register[2][4] ) );
  DLH_X1 \bank_register_reg[2][3]  ( .G(n3137), .D(n3152), .Q(
        \bank_register[2][3] ) );
  DLH_X1 \bank_register_reg[2][2]  ( .G(n3137), .D(n3149), .Q(
        \bank_register[2][2] ) );
  DLH_X1 \bank_register_reg[2][1]  ( .G(n3137), .D(n3146), .Q(
        \bank_register[2][1] ) );
  DLH_X1 \bank_register_reg[2][0]  ( .G(n3136), .D(n3143), .Q(
        \bank_register[2][0] ) );
  DLH_X1 \bank_register_reg[3][31]  ( .G(n3135), .D(n3236), .Q(
        \bank_register[3][31] ) );
  DLH_X1 \bank_register_reg[3][30]  ( .G(n3135), .D(n3233), .Q(
        \bank_register[3][30] ) );
  DLH_X1 \bank_register_reg[3][29]  ( .G(n3133), .D(n3230), .Q(
        \bank_register[3][29] ) );
  DLH_X1 \bank_register_reg[3][28]  ( .G(n3133), .D(n3227), .Q(
        \bank_register[3][28] ) );
  DLH_X1 \bank_register_reg[3][27]  ( .G(n3133), .D(n3224), .Q(
        \bank_register[3][27] ) );
  DLH_X1 \bank_register_reg[3][26]  ( .G(n3133), .D(n3221), .Q(
        \bank_register[3][26] ) );
  DLH_X1 \bank_register_reg[3][25]  ( .G(n3133), .D(n3218), .Q(
        \bank_register[3][25] ) );
  DLH_X1 \bank_register_reg[3][24]  ( .G(n3133), .D(n3215), .Q(
        \bank_register[3][24] ) );
  DLH_X1 \bank_register_reg[3][23]  ( .G(n3133), .D(n3212), .Q(
        \bank_register[3][23] ) );
  DLH_X1 \bank_register_reg[3][22]  ( .G(n3133), .D(n3209), .Q(
        \bank_register[3][22] ) );
  DLH_X1 \bank_register_reg[3][21]  ( .G(n3133), .D(n3206), .Q(
        \bank_register[3][21] ) );
  DLH_X1 \bank_register_reg[3][20]  ( .G(n3133), .D(n3203), .Q(
        \bank_register[3][20] ) );
  DLH_X1 \bank_register_reg[3][19]  ( .G(n3134), .D(n3200), .Q(
        \bank_register[3][19] ) );
  DLH_X1 \bank_register_reg[3][18]  ( .G(n3134), .D(n3197), .Q(
        \bank_register[3][18] ) );
  DLH_X1 \bank_register_reg[3][17]  ( .G(n3135), .D(n3194), .Q(
        \bank_register[3][17] ) );
  DLH_X1 \bank_register_reg[3][16]  ( .G(n3135), .D(n3191), .Q(
        \bank_register[3][16] ) );
  DLH_X1 \bank_register_reg[3][15]  ( .G(n3135), .D(n3188), .Q(
        \bank_register[3][15] ) );
  DLH_X1 \bank_register_reg[3][14]  ( .G(n3135), .D(n3185), .Q(
        \bank_register[3][14] ) );
  DLH_X1 \bank_register_reg[3][13]  ( .G(n3135), .D(n3182), .Q(
        \bank_register[3][13] ) );
  DLH_X1 \bank_register_reg[3][12]  ( .G(n3135), .D(n3179), .Q(
        \bank_register[3][12] ) );
  DLH_X1 \bank_register_reg[3][11]  ( .G(n3135), .D(n3176), .Q(
        \bank_register[3][11] ) );
  DLH_X1 \bank_register_reg[3][10]  ( .G(n3135), .D(n3173), .Q(
        \bank_register[3][10] ) );
  DLH_X1 \bank_register_reg[3][9]  ( .G(n3134), .D(n3170), .Q(
        \bank_register[3][9] ) );
  DLH_X1 \bank_register_reg[3][8]  ( .G(n3134), .D(n3167), .Q(
        \bank_register[3][8] ) );
  DLH_X1 \bank_register_reg[3][7]  ( .G(n3134), .D(n3164), .Q(
        \bank_register[3][7] ) );
  DLH_X1 \bank_register_reg[3][6]  ( .G(n3134), .D(n3161), .Q(
        \bank_register[3][6] ) );
  DLH_X1 \bank_register_reg[3][5]  ( .G(n3134), .D(n3158), .Q(
        \bank_register[3][5] ) );
  DLH_X1 \bank_register_reg[3][4]  ( .G(n3134), .D(n3155), .Q(
        \bank_register[3][4] ) );
  DLH_X1 \bank_register_reg[3][3]  ( .G(n3134), .D(n3152), .Q(
        \bank_register[3][3] ) );
  DLH_X1 \bank_register_reg[3][2]  ( .G(n3134), .D(n3149), .Q(
        \bank_register[3][2] ) );
  DLH_X1 \bank_register_reg[3][1]  ( .G(n3134), .D(n3146), .Q(
        \bank_register[3][1] ) );
  DLH_X1 \bank_register_reg[3][0]  ( .G(n3133), .D(n3143), .Q(
        \bank_register[3][0] ) );
  DLH_X1 \bank_register_reg[4][31]  ( .G(n3132), .D(n3236), .Q(
        \bank_register[4][31] ) );
  DLH_X1 \bank_register_reg[4][30]  ( .G(n3132), .D(n3233), .Q(
        \bank_register[4][30] ) );
  DLH_X1 \bank_register_reg[4][29]  ( .G(n3130), .D(n3230), .Q(
        \bank_register[4][29] ) );
  DLH_X1 \bank_register_reg[4][28]  ( .G(n3130), .D(n3227), .Q(
        \bank_register[4][28] ) );
  DLH_X1 \bank_register_reg[4][27]  ( .G(n3130), .D(n3224), .Q(
        \bank_register[4][27] ) );
  DLH_X1 \bank_register_reg[4][26]  ( .G(n3130), .D(n3221), .Q(
        \bank_register[4][26] ) );
  DLH_X1 \bank_register_reg[4][25]  ( .G(n3130), .D(n3218), .Q(
        \bank_register[4][25] ) );
  DLH_X1 \bank_register_reg[4][24]  ( .G(n3130), .D(n3215), .Q(
        \bank_register[4][24] ) );
  DLH_X1 \bank_register_reg[4][23]  ( .G(n3130), .D(n3212), .Q(
        \bank_register[4][23] ) );
  DLH_X1 \bank_register_reg[4][22]  ( .G(n3130), .D(n3209), .Q(
        \bank_register[4][22] ) );
  DLH_X1 \bank_register_reg[4][21]  ( .G(n3130), .D(n3206), .Q(
        \bank_register[4][21] ) );
  DLH_X1 \bank_register_reg[4][20]  ( .G(n3130), .D(n3203), .Q(
        \bank_register[4][20] ) );
  DLH_X1 \bank_register_reg[4][19]  ( .G(n3131), .D(n3200), .Q(
        \bank_register[4][19] ) );
  DLH_X1 \bank_register_reg[4][18]  ( .G(n3131), .D(n3197), .Q(
        \bank_register[4][18] ) );
  DLH_X1 \bank_register_reg[4][17]  ( .G(n3132), .D(n3194), .Q(
        \bank_register[4][17] ) );
  DLH_X1 \bank_register_reg[4][16]  ( .G(n3132), .D(n3191), .Q(
        \bank_register[4][16] ) );
  DLH_X1 \bank_register_reg[4][15]  ( .G(n3132), .D(n3188), .Q(
        \bank_register[4][15] ) );
  DLH_X1 \bank_register_reg[4][14]  ( .G(n3132), .D(n3185), .Q(
        \bank_register[4][14] ) );
  DLH_X1 \bank_register_reg[4][13]  ( .G(n3132), .D(n3182), .Q(
        \bank_register[4][13] ) );
  DLH_X1 \bank_register_reg[4][12]  ( .G(n3132), .D(n3179), .Q(
        \bank_register[4][12] ) );
  DLH_X1 \bank_register_reg[4][11]  ( .G(n3132), .D(n3176), .Q(
        \bank_register[4][11] ) );
  DLH_X1 \bank_register_reg[4][10]  ( .G(n3132), .D(n3173), .Q(
        \bank_register[4][10] ) );
  DLH_X1 \bank_register_reg[4][9]  ( .G(n3131), .D(n3170), .Q(
        \bank_register[4][9] ) );
  DLH_X1 \bank_register_reg[4][8]  ( .G(n3131), .D(n3167), .Q(
        \bank_register[4][8] ) );
  DLH_X1 \bank_register_reg[4][7]  ( .G(n3131), .D(n3164), .Q(
        \bank_register[4][7] ) );
  DLH_X1 \bank_register_reg[4][6]  ( .G(n3131), .D(n3161), .Q(
        \bank_register[4][6] ) );
  DLH_X1 \bank_register_reg[4][5]  ( .G(n3131), .D(n3158), .Q(
        \bank_register[4][5] ) );
  DLH_X1 \bank_register_reg[4][4]  ( .G(n3131), .D(n3155), .Q(
        \bank_register[4][4] ) );
  DLH_X1 \bank_register_reg[4][3]  ( .G(n3131), .D(n3152), .Q(
        \bank_register[4][3] ) );
  DLH_X1 \bank_register_reg[4][2]  ( .G(n3131), .D(n3149), .Q(
        \bank_register[4][2] ) );
  DLH_X1 \bank_register_reg[4][1]  ( .G(n3131), .D(n3146), .Q(
        \bank_register[4][1] ) );
  DLH_X1 \bank_register_reg[4][0]  ( .G(n3130), .D(n3143), .Q(
        \bank_register[4][0] ) );
  DLH_X1 \bank_register_reg[5][31]  ( .G(n3129), .D(n3236), .Q(
        \bank_register[5][31] ) );
  DLH_X1 \bank_register_reg[5][30]  ( .G(n3129), .D(n3233), .Q(
        \bank_register[5][30] ) );
  DLH_X1 \bank_register_reg[5][29]  ( .G(n3127), .D(n3230), .Q(
        \bank_register[5][29] ) );
  DLH_X1 \bank_register_reg[5][28]  ( .G(n3127), .D(n3227), .Q(
        \bank_register[5][28] ) );
  DLH_X1 \bank_register_reg[5][27]  ( .G(n3127), .D(n3224), .Q(
        \bank_register[5][27] ) );
  DLH_X1 \bank_register_reg[5][26]  ( .G(n3127), .D(n3221), .Q(
        \bank_register[5][26] ) );
  DLH_X1 \bank_register_reg[5][25]  ( .G(n3127), .D(n3218), .Q(
        \bank_register[5][25] ) );
  DLH_X1 \bank_register_reg[5][24]  ( .G(n3127), .D(n3215), .Q(
        \bank_register[5][24] ) );
  DLH_X1 \bank_register_reg[5][23]  ( .G(n3127), .D(n3212), .Q(
        \bank_register[5][23] ) );
  DLH_X1 \bank_register_reg[5][22]  ( .G(n3127), .D(n3209), .Q(
        \bank_register[5][22] ) );
  DLH_X1 \bank_register_reg[5][21]  ( .G(n3127), .D(n3206), .Q(
        \bank_register[5][21] ) );
  DLH_X1 \bank_register_reg[5][20]  ( .G(n3127), .D(n3203), .Q(
        \bank_register[5][20] ) );
  DLH_X1 \bank_register_reg[5][19]  ( .G(n3128), .D(n3200), .Q(
        \bank_register[5][19] ) );
  DLH_X1 \bank_register_reg[5][18]  ( .G(n3128), .D(n3197), .Q(
        \bank_register[5][18] ) );
  DLH_X1 \bank_register_reg[5][17]  ( .G(n3129), .D(n3194), .Q(
        \bank_register[5][17] ) );
  DLH_X1 \bank_register_reg[5][16]  ( .G(n3129), .D(n3191), .Q(
        \bank_register[5][16] ) );
  DLH_X1 \bank_register_reg[5][15]  ( .G(n3129), .D(n3188), .Q(
        \bank_register[5][15] ) );
  DLH_X1 \bank_register_reg[5][14]  ( .G(n3129), .D(n3185), .Q(
        \bank_register[5][14] ) );
  DLH_X1 \bank_register_reg[5][13]  ( .G(n3129), .D(n3182), .Q(
        \bank_register[5][13] ) );
  DLH_X1 \bank_register_reg[5][12]  ( .G(n3129), .D(n3179), .Q(
        \bank_register[5][12] ) );
  DLH_X1 \bank_register_reg[5][11]  ( .G(n3129), .D(n3176), .Q(
        \bank_register[5][11] ) );
  DLH_X1 \bank_register_reg[5][10]  ( .G(n3129), .D(n3173), .Q(
        \bank_register[5][10] ) );
  DLH_X1 \bank_register_reg[5][9]  ( .G(n3128), .D(n3170), .Q(
        \bank_register[5][9] ) );
  DLH_X1 \bank_register_reg[5][8]  ( .G(n3128), .D(n3167), .Q(
        \bank_register[5][8] ) );
  DLH_X1 \bank_register_reg[5][7]  ( .G(n3128), .D(n3164), .Q(
        \bank_register[5][7] ) );
  DLH_X1 \bank_register_reg[5][6]  ( .G(n3128), .D(n3161), .Q(
        \bank_register[5][6] ) );
  DLH_X1 \bank_register_reg[5][5]  ( .G(n3128), .D(n3158), .Q(
        \bank_register[5][5] ) );
  DLH_X1 \bank_register_reg[5][4]  ( .G(n3128), .D(n3155), .Q(
        \bank_register[5][4] ) );
  DLH_X1 \bank_register_reg[5][3]  ( .G(n3128), .D(n3152), .Q(
        \bank_register[5][3] ) );
  DLH_X1 \bank_register_reg[5][2]  ( .G(n3128), .D(n3149), .Q(
        \bank_register[5][2] ) );
  DLH_X1 \bank_register_reg[5][1]  ( .G(n3128), .D(n3146), .Q(
        \bank_register[5][1] ) );
  DLH_X1 \bank_register_reg[5][0]  ( .G(n3127), .D(n3143), .Q(
        \bank_register[5][0] ) );
  DLH_X1 \bank_register_reg[6][31]  ( .G(n3126), .D(n3236), .Q(
        \bank_register[6][31] ) );
  DLH_X1 \bank_register_reg[6][30]  ( .G(n3126), .D(n3233), .Q(
        \bank_register[6][30] ) );
  DLH_X1 \bank_register_reg[6][29]  ( .G(n3124), .D(n3230), .Q(
        \bank_register[6][29] ) );
  DLH_X1 \bank_register_reg[6][28]  ( .G(n3124), .D(n3227), .Q(
        \bank_register[6][28] ) );
  DLH_X1 \bank_register_reg[6][27]  ( .G(n3124), .D(n3224), .Q(
        \bank_register[6][27] ) );
  DLH_X1 \bank_register_reg[6][26]  ( .G(n3124), .D(n3221), .Q(
        \bank_register[6][26] ) );
  DLH_X1 \bank_register_reg[6][25]  ( .G(n3124), .D(n3218), .Q(
        \bank_register[6][25] ) );
  DLH_X1 \bank_register_reg[6][24]  ( .G(n3124), .D(n3215), .Q(
        \bank_register[6][24] ) );
  DLH_X1 \bank_register_reg[6][23]  ( .G(n3124), .D(n3212), .Q(
        \bank_register[6][23] ) );
  DLH_X1 \bank_register_reg[6][22]  ( .G(n3124), .D(n3209), .Q(
        \bank_register[6][22] ) );
  DLH_X1 \bank_register_reg[6][21]  ( .G(n3124), .D(n3206), .Q(
        \bank_register[6][21] ) );
  DLH_X1 \bank_register_reg[6][20]  ( .G(n3124), .D(n3203), .Q(
        \bank_register[6][20] ) );
  DLH_X1 \bank_register_reg[6][19]  ( .G(n3125), .D(n3200), .Q(
        \bank_register[6][19] ) );
  DLH_X1 \bank_register_reg[6][18]  ( .G(n3125), .D(n3197), .Q(
        \bank_register[6][18] ) );
  DLH_X1 \bank_register_reg[6][17]  ( .G(n3126), .D(n3194), .Q(
        \bank_register[6][17] ) );
  DLH_X1 \bank_register_reg[6][16]  ( .G(n3126), .D(n3191), .Q(
        \bank_register[6][16] ) );
  DLH_X1 \bank_register_reg[6][15]  ( .G(n3126), .D(n3188), .Q(
        \bank_register[6][15] ) );
  DLH_X1 \bank_register_reg[6][14]  ( .G(n3126), .D(n3185), .Q(
        \bank_register[6][14] ) );
  DLH_X1 \bank_register_reg[6][13]  ( .G(n3126), .D(n3182), .Q(
        \bank_register[6][13] ) );
  DLH_X1 \bank_register_reg[6][12]  ( .G(n3126), .D(n3179), .Q(
        \bank_register[6][12] ) );
  DLH_X1 \bank_register_reg[6][11]  ( .G(n3126), .D(n3176), .Q(
        \bank_register[6][11] ) );
  DLH_X1 \bank_register_reg[6][10]  ( .G(n3126), .D(n3173), .Q(
        \bank_register[6][10] ) );
  DLH_X1 \bank_register_reg[6][9]  ( .G(n3125), .D(n3170), .Q(
        \bank_register[6][9] ) );
  DLH_X1 \bank_register_reg[6][8]  ( .G(n3125), .D(n3167), .Q(
        \bank_register[6][8] ) );
  DLH_X1 \bank_register_reg[6][7]  ( .G(n3125), .D(n3164), .Q(
        \bank_register[6][7] ) );
  DLH_X1 \bank_register_reg[6][6]  ( .G(n3125), .D(n3161), .Q(
        \bank_register[6][6] ) );
  DLH_X1 \bank_register_reg[6][5]  ( .G(n3125), .D(n3158), .Q(
        \bank_register[6][5] ) );
  DLH_X1 \bank_register_reg[6][4]  ( .G(n3125), .D(n3155), .Q(
        \bank_register[6][4] ) );
  DLH_X1 \bank_register_reg[6][3]  ( .G(n3125), .D(n3152), .Q(
        \bank_register[6][3] ) );
  DLH_X1 \bank_register_reg[6][2]  ( .G(n3125), .D(n3149), .Q(
        \bank_register[6][2] ) );
  DLH_X1 \bank_register_reg[6][1]  ( .G(n3125), .D(n3146), .Q(
        \bank_register[6][1] ) );
  DLH_X1 \bank_register_reg[6][0]  ( .G(n3124), .D(n3143), .Q(
        \bank_register[6][0] ) );
  DLH_X1 \bank_register_reg[7][31]  ( .G(n3123), .D(n3236), .Q(
        \bank_register[7][31] ) );
  DLH_X1 \bank_register_reg[7][30]  ( .G(n3123), .D(n3233), .Q(
        \bank_register[7][30] ) );
  DLH_X1 \bank_register_reg[7][29]  ( .G(n3121), .D(n3230), .Q(
        \bank_register[7][29] ) );
  DLH_X1 \bank_register_reg[7][28]  ( .G(n3121), .D(n3227), .Q(
        \bank_register[7][28] ) );
  DLH_X1 \bank_register_reg[7][27]  ( .G(n3121), .D(n3224), .Q(
        \bank_register[7][27] ) );
  DLH_X1 \bank_register_reg[7][26]  ( .G(n3121), .D(n3221), .Q(
        \bank_register[7][26] ) );
  DLH_X1 \bank_register_reg[7][25]  ( .G(n3121), .D(n3218), .Q(
        \bank_register[7][25] ) );
  DLH_X1 \bank_register_reg[7][24]  ( .G(n3121), .D(n3215), .Q(
        \bank_register[7][24] ) );
  DLH_X1 \bank_register_reg[7][23]  ( .G(n3121), .D(n3212), .Q(
        \bank_register[7][23] ) );
  DLH_X1 \bank_register_reg[7][22]  ( .G(n3121), .D(n3209), .Q(
        \bank_register[7][22] ) );
  DLH_X1 \bank_register_reg[7][21]  ( .G(n3121), .D(n3206), .Q(
        \bank_register[7][21] ) );
  DLH_X1 \bank_register_reg[7][20]  ( .G(n3121), .D(n3203), .Q(
        \bank_register[7][20] ) );
  DLH_X1 \bank_register_reg[7][19]  ( .G(n3122), .D(n3200), .Q(
        \bank_register[7][19] ) );
  DLH_X1 \bank_register_reg[7][18]  ( .G(n3122), .D(n3197), .Q(
        \bank_register[7][18] ) );
  DLH_X1 \bank_register_reg[7][17]  ( .G(n3123), .D(n3194), .Q(
        \bank_register[7][17] ) );
  DLH_X1 \bank_register_reg[7][16]  ( .G(n3123), .D(n3191), .Q(
        \bank_register[7][16] ) );
  DLH_X1 \bank_register_reg[7][15]  ( .G(n3123), .D(n3188), .Q(
        \bank_register[7][15] ) );
  DLH_X1 \bank_register_reg[7][14]  ( .G(n3123), .D(n3185), .Q(
        \bank_register[7][14] ) );
  DLH_X1 \bank_register_reg[7][13]  ( .G(n3123), .D(n3182), .Q(
        \bank_register[7][13] ) );
  DLH_X1 \bank_register_reg[7][12]  ( .G(n3123), .D(n3179), .Q(
        \bank_register[7][12] ) );
  DLH_X1 \bank_register_reg[7][11]  ( .G(n3123), .D(n3176), .Q(
        \bank_register[7][11] ) );
  DLH_X1 \bank_register_reg[7][10]  ( .G(n3123), .D(n3173), .Q(
        \bank_register[7][10] ) );
  DLH_X1 \bank_register_reg[7][9]  ( .G(n3122), .D(n3170), .Q(
        \bank_register[7][9] ) );
  DLH_X1 \bank_register_reg[7][8]  ( .G(n3122), .D(n3167), .Q(
        \bank_register[7][8] ) );
  DLH_X1 \bank_register_reg[7][7]  ( .G(n3122), .D(n3164), .Q(
        \bank_register[7][7] ) );
  DLH_X1 \bank_register_reg[7][6]  ( .G(n3122), .D(n3161), .Q(
        \bank_register[7][6] ) );
  DLH_X1 \bank_register_reg[7][5]  ( .G(n3122), .D(n3158), .Q(
        \bank_register[7][5] ) );
  DLH_X1 \bank_register_reg[7][4]  ( .G(n3122), .D(n3155), .Q(
        \bank_register[7][4] ) );
  DLH_X1 \bank_register_reg[7][3]  ( .G(n3122), .D(n3152), .Q(
        \bank_register[7][3] ) );
  DLH_X1 \bank_register_reg[7][2]  ( .G(n3122), .D(n3149), .Q(
        \bank_register[7][2] ) );
  DLH_X1 \bank_register_reg[7][1]  ( .G(n3122), .D(n3146), .Q(
        \bank_register[7][1] ) );
  DLH_X1 \bank_register_reg[7][0]  ( .G(n3121), .D(n3143), .Q(
        \bank_register[7][0] ) );
  DLH_X1 \bank_register_reg[8][31]  ( .G(n3120), .D(n3236), .Q(
        \bank_register[8][31] ) );
  DLH_X1 \bank_register_reg[8][30]  ( .G(n3120), .D(n3233), .Q(
        \bank_register[8][30] ) );
  DLH_X1 \bank_register_reg[8][29]  ( .G(n3118), .D(n3230), .Q(
        \bank_register[8][29] ) );
  DLH_X1 \bank_register_reg[8][28]  ( .G(n3118), .D(n3227), .Q(
        \bank_register[8][28] ) );
  DLH_X1 \bank_register_reg[8][27]  ( .G(n3118), .D(n3224), .Q(
        \bank_register[8][27] ) );
  DLH_X1 \bank_register_reg[8][26]  ( .G(n3118), .D(n3221), .Q(
        \bank_register[8][26] ) );
  DLH_X1 \bank_register_reg[8][25]  ( .G(n3118), .D(n3218), .Q(
        \bank_register[8][25] ) );
  DLH_X1 \bank_register_reg[8][24]  ( .G(n3118), .D(n3215), .Q(
        \bank_register[8][24] ) );
  DLH_X1 \bank_register_reg[8][23]  ( .G(n3118), .D(n3212), .Q(
        \bank_register[8][23] ) );
  DLH_X1 \bank_register_reg[8][22]  ( .G(n3118), .D(n3209), .Q(
        \bank_register[8][22] ) );
  DLH_X1 \bank_register_reg[8][21]  ( .G(n3118), .D(n3206), .Q(
        \bank_register[8][21] ) );
  DLH_X1 \bank_register_reg[8][20]  ( .G(n3118), .D(n3203), .Q(
        \bank_register[8][20] ) );
  DLH_X1 \bank_register_reg[8][19]  ( .G(n3119), .D(n3200), .Q(
        \bank_register[8][19] ) );
  DLH_X1 \bank_register_reg[8][18]  ( .G(n3119), .D(n3197), .Q(
        \bank_register[8][18] ) );
  DLH_X1 \bank_register_reg[8][17]  ( .G(n3120), .D(n3194), .Q(
        \bank_register[8][17] ) );
  DLH_X1 \bank_register_reg[8][16]  ( .G(n3120), .D(n3191), .Q(
        \bank_register[8][16] ) );
  DLH_X1 \bank_register_reg[8][15]  ( .G(n3120), .D(n3188), .Q(
        \bank_register[8][15] ) );
  DLH_X1 \bank_register_reg[8][14]  ( .G(n3120), .D(n3185), .Q(
        \bank_register[8][14] ) );
  DLH_X1 \bank_register_reg[8][13]  ( .G(n3120), .D(n3182), .Q(
        \bank_register[8][13] ) );
  DLH_X1 \bank_register_reg[8][12]  ( .G(n3120), .D(n3179), .Q(
        \bank_register[8][12] ) );
  DLH_X1 \bank_register_reg[8][11]  ( .G(n3120), .D(n3176), .Q(
        \bank_register[8][11] ) );
  DLH_X1 \bank_register_reg[8][10]  ( .G(n3120), .D(n3173), .Q(
        \bank_register[8][10] ) );
  DLH_X1 \bank_register_reg[8][9]  ( .G(n3119), .D(n3170), .Q(
        \bank_register[8][9] ) );
  DLH_X1 \bank_register_reg[8][8]  ( .G(n3119), .D(n3167), .Q(
        \bank_register[8][8] ) );
  DLH_X1 \bank_register_reg[8][7]  ( .G(n3119), .D(n3164), .Q(
        \bank_register[8][7] ) );
  DLH_X1 \bank_register_reg[8][6]  ( .G(n3119), .D(n3161), .Q(
        \bank_register[8][6] ) );
  DLH_X1 \bank_register_reg[8][5]  ( .G(n3119), .D(n3158), .Q(
        \bank_register[8][5] ) );
  DLH_X1 \bank_register_reg[8][4]  ( .G(n3119), .D(n3155), .Q(
        \bank_register[8][4] ) );
  DLH_X1 \bank_register_reg[8][3]  ( .G(n3119), .D(n3152), .Q(
        \bank_register[8][3] ) );
  DLH_X1 \bank_register_reg[8][2]  ( .G(n3119), .D(n3149), .Q(
        \bank_register[8][2] ) );
  DLH_X1 \bank_register_reg[8][1]  ( .G(n3119), .D(n3146), .Q(
        \bank_register[8][1] ) );
  DLH_X1 \bank_register_reg[8][0]  ( .G(n3118), .D(n3143), .Q(
        \bank_register[8][0] ) );
  DLH_X1 \bank_register_reg[9][31]  ( .G(n3117), .D(n3236), .Q(
        \bank_register[9][31] ) );
  DLH_X1 \bank_register_reg[9][30]  ( .G(n3117), .D(n3233), .Q(
        \bank_register[9][30] ) );
  DLH_X1 \bank_register_reg[9][29]  ( .G(n3115), .D(n3230), .Q(
        \bank_register[9][29] ) );
  DLH_X1 \bank_register_reg[9][28]  ( .G(n3115), .D(n3227), .Q(
        \bank_register[9][28] ) );
  DLH_X1 \bank_register_reg[9][27]  ( .G(n3115), .D(n3224), .Q(
        \bank_register[9][27] ) );
  DLH_X1 \bank_register_reg[9][26]  ( .G(n3115), .D(n3221), .Q(
        \bank_register[9][26] ) );
  DLH_X1 \bank_register_reg[9][25]  ( .G(n3115), .D(n3218), .Q(
        \bank_register[9][25] ) );
  DLH_X1 \bank_register_reg[9][24]  ( .G(n3115), .D(n3215), .Q(
        \bank_register[9][24] ) );
  DLH_X1 \bank_register_reg[9][23]  ( .G(n3115), .D(n3212), .Q(
        \bank_register[9][23] ) );
  DLH_X1 \bank_register_reg[9][22]  ( .G(n3115), .D(n3209), .Q(
        \bank_register[9][22] ) );
  DLH_X1 \bank_register_reg[9][21]  ( .G(n3115), .D(n3206), .Q(
        \bank_register[9][21] ) );
  DLH_X1 \bank_register_reg[9][20]  ( .G(n3115), .D(n3203), .Q(
        \bank_register[9][20] ) );
  DLH_X1 \bank_register_reg[9][19]  ( .G(n3116), .D(n3200), .Q(
        \bank_register[9][19] ) );
  DLH_X1 \bank_register_reg[9][18]  ( .G(n3116), .D(n3197), .Q(
        \bank_register[9][18] ) );
  DLH_X1 \bank_register_reg[9][17]  ( .G(n3117), .D(n3194), .Q(
        \bank_register[9][17] ) );
  DLH_X1 \bank_register_reg[9][16]  ( .G(n3117), .D(n3191), .Q(
        \bank_register[9][16] ) );
  DLH_X1 \bank_register_reg[9][15]  ( .G(n3117), .D(n3188), .Q(
        \bank_register[9][15] ) );
  DLH_X1 \bank_register_reg[9][14]  ( .G(n3117), .D(n3185), .Q(
        \bank_register[9][14] ) );
  DLH_X1 \bank_register_reg[9][13]  ( .G(n3117), .D(n3182), .Q(
        \bank_register[9][13] ) );
  DLH_X1 \bank_register_reg[9][12]  ( .G(n3117), .D(n3179), .Q(
        \bank_register[9][12] ) );
  DLH_X1 \bank_register_reg[9][11]  ( .G(n3117), .D(n3176), .Q(
        \bank_register[9][11] ) );
  DLH_X1 \bank_register_reg[9][10]  ( .G(n3117), .D(n3173), .Q(
        \bank_register[9][10] ) );
  DLH_X1 \bank_register_reg[9][9]  ( .G(n3116), .D(n3170), .Q(
        \bank_register[9][9] ) );
  DLH_X1 \bank_register_reg[9][8]  ( .G(n3116), .D(n3167), .Q(
        \bank_register[9][8] ) );
  DLH_X1 \bank_register_reg[9][7]  ( .G(n3116), .D(n3164), .Q(
        \bank_register[9][7] ) );
  DLH_X1 \bank_register_reg[9][6]  ( .G(n3116), .D(n3161), .Q(
        \bank_register[9][6] ) );
  DLH_X1 \bank_register_reg[9][5]  ( .G(n3116), .D(n3158), .Q(
        \bank_register[9][5] ) );
  DLH_X1 \bank_register_reg[9][4]  ( .G(n3116), .D(n3155), .Q(
        \bank_register[9][4] ) );
  DLH_X1 \bank_register_reg[9][3]  ( .G(n3116), .D(n3152), .Q(
        \bank_register[9][3] ) );
  DLH_X1 \bank_register_reg[9][2]  ( .G(n3116), .D(n3149), .Q(
        \bank_register[9][2] ) );
  DLH_X1 \bank_register_reg[9][1]  ( .G(n3116), .D(n3146), .Q(
        \bank_register[9][1] ) );
  DLH_X1 \bank_register_reg[9][0]  ( .G(n3115), .D(n3143), .Q(
        \bank_register[9][0] ) );
  DLH_X1 \bank_register_reg[10][31]  ( .G(n3114), .D(n3236), .Q(
        \bank_register[10][31] ) );
  DLH_X1 \bank_register_reg[10][30]  ( .G(n3114), .D(n3233), .Q(
        \bank_register[10][30] ) );
  DLH_X1 \bank_register_reg[10][29]  ( .G(n3112), .D(n3230), .Q(
        \bank_register[10][29] ) );
  DLH_X1 \bank_register_reg[10][28]  ( .G(n3112), .D(n3227), .Q(
        \bank_register[10][28] ) );
  DLH_X1 \bank_register_reg[10][27]  ( .G(n3112), .D(n3224), .Q(
        \bank_register[10][27] ) );
  DLH_X1 \bank_register_reg[10][26]  ( .G(n3112), .D(n3221), .Q(
        \bank_register[10][26] ) );
  DLH_X1 \bank_register_reg[10][25]  ( .G(n3112), .D(n3218), .Q(
        \bank_register[10][25] ) );
  DLH_X1 \bank_register_reg[10][24]  ( .G(n3112), .D(n3215), .Q(
        \bank_register[10][24] ) );
  DLH_X1 \bank_register_reg[10][23]  ( .G(n3112), .D(n3212), .Q(
        \bank_register[10][23] ) );
  DLH_X1 \bank_register_reg[10][22]  ( .G(n3112), .D(n3209), .Q(
        \bank_register[10][22] ) );
  DLH_X1 \bank_register_reg[10][21]  ( .G(n3112), .D(n3206), .Q(
        \bank_register[10][21] ) );
  DLH_X1 \bank_register_reg[10][20]  ( .G(n3112), .D(n3203), .Q(
        \bank_register[10][20] ) );
  DLH_X1 \bank_register_reg[10][19]  ( .G(n3113), .D(n3200), .Q(
        \bank_register[10][19] ) );
  DLH_X1 \bank_register_reg[10][18]  ( .G(n3113), .D(n3197), .Q(
        \bank_register[10][18] ) );
  DLH_X1 \bank_register_reg[10][17]  ( .G(n3114), .D(n3194), .Q(
        \bank_register[10][17] ) );
  DLH_X1 \bank_register_reg[10][16]  ( .G(n3114), .D(n3191), .Q(
        \bank_register[10][16] ) );
  DLH_X1 \bank_register_reg[10][15]  ( .G(n3114), .D(n3188), .Q(
        \bank_register[10][15] ) );
  DLH_X1 \bank_register_reg[10][14]  ( .G(n3114), .D(n3185), .Q(
        \bank_register[10][14] ) );
  DLH_X1 \bank_register_reg[10][13]  ( .G(n3114), .D(n3182), .Q(
        \bank_register[10][13] ) );
  DLH_X1 \bank_register_reg[10][12]  ( .G(n3114), .D(n3179), .Q(
        \bank_register[10][12] ) );
  DLH_X1 \bank_register_reg[10][11]  ( .G(n3114), .D(n3176), .Q(
        \bank_register[10][11] ) );
  DLH_X1 \bank_register_reg[10][10]  ( .G(n3114), .D(n3173), .Q(
        \bank_register[10][10] ) );
  DLH_X1 \bank_register_reg[10][9]  ( .G(n3113), .D(n3170), .Q(
        \bank_register[10][9] ) );
  DLH_X1 \bank_register_reg[10][8]  ( .G(n3113), .D(n3167), .Q(
        \bank_register[10][8] ) );
  DLH_X1 \bank_register_reg[10][7]  ( .G(n3113), .D(n3164), .Q(
        \bank_register[10][7] ) );
  DLH_X1 \bank_register_reg[10][6]  ( .G(n3113), .D(n3161), .Q(
        \bank_register[10][6] ) );
  DLH_X1 \bank_register_reg[10][5]  ( .G(n3113), .D(n3158), .Q(
        \bank_register[10][5] ) );
  DLH_X1 \bank_register_reg[10][4]  ( .G(n3113), .D(n3155), .Q(
        \bank_register[10][4] ) );
  DLH_X1 \bank_register_reg[10][3]  ( .G(n3113), .D(n3152), .Q(
        \bank_register[10][3] ) );
  DLH_X1 \bank_register_reg[10][2]  ( .G(n3113), .D(n3149), .Q(
        \bank_register[10][2] ) );
  DLH_X1 \bank_register_reg[10][1]  ( .G(n3113), .D(n3146), .Q(
        \bank_register[10][1] ) );
  DLH_X1 \bank_register_reg[10][0]  ( .G(n3112), .D(n3143), .Q(
        \bank_register[10][0] ) );
  DLH_X1 \bank_register_reg[11][31]  ( .G(n3111), .D(n3237), .Q(
        \bank_register[11][31] ) );
  DLH_X1 \bank_register_reg[11][30]  ( .G(n3111), .D(n3234), .Q(
        \bank_register[11][30] ) );
  DLH_X1 \bank_register_reg[11][29]  ( .G(n3109), .D(n3231), .Q(
        \bank_register[11][29] ) );
  DLH_X1 \bank_register_reg[11][28]  ( .G(n3109), .D(n3228), .Q(
        \bank_register[11][28] ) );
  DLH_X1 \bank_register_reg[11][27]  ( .G(n3109), .D(n3225), .Q(
        \bank_register[11][27] ) );
  DLH_X1 \bank_register_reg[11][26]  ( .G(n3109), .D(n3222), .Q(
        \bank_register[11][26] ) );
  DLH_X1 \bank_register_reg[11][25]  ( .G(n3109), .D(n3219), .Q(
        \bank_register[11][25] ) );
  DLH_X1 \bank_register_reg[11][24]  ( .G(n3109), .D(n3216), .Q(
        \bank_register[11][24] ) );
  DLH_X1 \bank_register_reg[11][23]  ( .G(n3109), .D(n3213), .Q(
        \bank_register[11][23] ) );
  DLH_X1 \bank_register_reg[11][22]  ( .G(n3109), .D(n3210), .Q(
        \bank_register[11][22] ) );
  DLH_X1 \bank_register_reg[11][21]  ( .G(n3109), .D(n3207), .Q(
        \bank_register[11][21] ) );
  DLH_X1 \bank_register_reg[11][20]  ( .G(n3109), .D(n3204), .Q(
        \bank_register[11][20] ) );
  DLH_X1 \bank_register_reg[11][19]  ( .G(n3110), .D(n3201), .Q(
        \bank_register[11][19] ) );
  DLH_X1 \bank_register_reg[11][18]  ( .G(n3110), .D(n3198), .Q(
        \bank_register[11][18] ) );
  DLH_X1 \bank_register_reg[11][17]  ( .G(n3111), .D(n3195), .Q(
        \bank_register[11][17] ) );
  DLH_X1 \bank_register_reg[11][16]  ( .G(n3111), .D(n3192), .Q(
        \bank_register[11][16] ) );
  DLH_X1 \bank_register_reg[11][15]  ( .G(n3111), .D(n3189), .Q(
        \bank_register[11][15] ) );
  DLH_X1 \bank_register_reg[11][14]  ( .G(n3111), .D(n3186), .Q(
        \bank_register[11][14] ) );
  DLH_X1 \bank_register_reg[11][13]  ( .G(n3111), .D(n3183), .Q(
        \bank_register[11][13] ) );
  DLH_X1 \bank_register_reg[11][12]  ( .G(n3111), .D(n3180), .Q(
        \bank_register[11][12] ) );
  DLH_X1 \bank_register_reg[11][11]  ( .G(n3111), .D(n3177), .Q(
        \bank_register[11][11] ) );
  DLH_X1 \bank_register_reg[11][10]  ( .G(n3111), .D(n3174), .Q(
        \bank_register[11][10] ) );
  DLH_X1 \bank_register_reg[11][9]  ( .G(n3110), .D(n3171), .Q(
        \bank_register[11][9] ) );
  DLH_X1 \bank_register_reg[11][8]  ( .G(n3110), .D(n3168), .Q(
        \bank_register[11][8] ) );
  DLH_X1 \bank_register_reg[11][7]  ( .G(n3110), .D(n3165), .Q(
        \bank_register[11][7] ) );
  DLH_X1 \bank_register_reg[11][6]  ( .G(n3110), .D(n3162), .Q(
        \bank_register[11][6] ) );
  DLH_X1 \bank_register_reg[11][5]  ( .G(n3110), .D(n3159), .Q(
        \bank_register[11][5] ) );
  DLH_X1 \bank_register_reg[11][4]  ( .G(n3110), .D(n3156), .Q(
        \bank_register[11][4] ) );
  DLH_X1 \bank_register_reg[11][3]  ( .G(n3110), .D(n3153), .Q(
        \bank_register[11][3] ) );
  DLH_X1 \bank_register_reg[11][2]  ( .G(n3110), .D(n3150), .Q(
        \bank_register[11][2] ) );
  DLH_X1 \bank_register_reg[11][1]  ( .G(n3110), .D(n3147), .Q(
        \bank_register[11][1] ) );
  DLH_X1 \bank_register_reg[11][0]  ( .G(n3109), .D(n3144), .Q(
        \bank_register[11][0] ) );
  DLH_X1 \bank_register_reg[12][31]  ( .G(n3108), .D(n3237), .Q(
        \bank_register[12][31] ) );
  DLH_X1 \bank_register_reg[12][30]  ( .G(n3108), .D(n3234), .Q(
        \bank_register[12][30] ) );
  DLH_X1 \bank_register_reg[12][29]  ( .G(n3106), .D(n3231), .Q(
        \bank_register[12][29] ) );
  DLH_X1 \bank_register_reg[12][28]  ( .G(n3106), .D(n3228), .Q(
        \bank_register[12][28] ) );
  DLH_X1 \bank_register_reg[12][27]  ( .G(n3106), .D(n3225), .Q(
        \bank_register[12][27] ) );
  DLH_X1 \bank_register_reg[12][26]  ( .G(n3106), .D(n3222), .Q(
        \bank_register[12][26] ) );
  DLH_X1 \bank_register_reg[12][25]  ( .G(n3106), .D(n3219), .Q(
        \bank_register[12][25] ) );
  DLH_X1 \bank_register_reg[12][24]  ( .G(n3106), .D(n3216), .Q(
        \bank_register[12][24] ) );
  DLH_X1 \bank_register_reg[12][23]  ( .G(n3106), .D(n3213), .Q(
        \bank_register[12][23] ) );
  DLH_X1 \bank_register_reg[12][22]  ( .G(n3106), .D(n3210), .Q(
        \bank_register[12][22] ) );
  DLH_X1 \bank_register_reg[12][21]  ( .G(n3106), .D(n3207), .Q(
        \bank_register[12][21] ) );
  DLH_X1 \bank_register_reg[12][20]  ( .G(n3106), .D(n3204), .Q(
        \bank_register[12][20] ) );
  DLH_X1 \bank_register_reg[12][19]  ( .G(n3107), .D(n3201), .Q(
        \bank_register[12][19] ) );
  DLH_X1 \bank_register_reg[12][18]  ( .G(n3107), .D(n3198), .Q(
        \bank_register[12][18] ) );
  DLH_X1 \bank_register_reg[12][17]  ( .G(n3108), .D(n3195), .Q(
        \bank_register[12][17] ) );
  DLH_X1 \bank_register_reg[12][16]  ( .G(n3108), .D(n3192), .Q(
        \bank_register[12][16] ) );
  DLH_X1 \bank_register_reg[12][15]  ( .G(n3108), .D(n3189), .Q(
        \bank_register[12][15] ) );
  DLH_X1 \bank_register_reg[12][14]  ( .G(n3108), .D(n3186), .Q(
        \bank_register[12][14] ) );
  DLH_X1 \bank_register_reg[12][13]  ( .G(n3108), .D(n3183), .Q(
        \bank_register[12][13] ) );
  DLH_X1 \bank_register_reg[12][12]  ( .G(n3108), .D(n3180), .Q(
        \bank_register[12][12] ) );
  DLH_X1 \bank_register_reg[12][11]  ( .G(n3108), .D(n3177), .Q(
        \bank_register[12][11] ) );
  DLH_X1 \bank_register_reg[12][10]  ( .G(n3108), .D(n3174), .Q(
        \bank_register[12][10] ) );
  DLH_X1 \bank_register_reg[12][9]  ( .G(n3107), .D(n3171), .Q(
        \bank_register[12][9] ) );
  DLH_X1 \bank_register_reg[12][8]  ( .G(n3107), .D(n3168), .Q(
        \bank_register[12][8] ) );
  DLH_X1 \bank_register_reg[12][7]  ( .G(n3107), .D(n3165), .Q(
        \bank_register[12][7] ) );
  DLH_X1 \bank_register_reg[12][6]  ( .G(n3107), .D(n3162), .Q(
        \bank_register[12][6] ) );
  DLH_X1 \bank_register_reg[12][5]  ( .G(n3107), .D(n3159), .Q(
        \bank_register[12][5] ) );
  DLH_X1 \bank_register_reg[12][4]  ( .G(n3107), .D(n3156), .Q(
        \bank_register[12][4] ) );
  DLH_X1 \bank_register_reg[12][3]  ( .G(n3107), .D(n3153), .Q(
        \bank_register[12][3] ) );
  DLH_X1 \bank_register_reg[12][2]  ( .G(n3107), .D(n3150), .Q(
        \bank_register[12][2] ) );
  DLH_X1 \bank_register_reg[12][1]  ( .G(n3107), .D(n3147), .Q(
        \bank_register[12][1] ) );
  DLH_X1 \bank_register_reg[12][0]  ( .G(n3106), .D(n3144), .Q(
        \bank_register[12][0] ) );
  DLH_X1 \bank_register_reg[13][31]  ( .G(n3105), .D(n3237), .Q(
        \bank_register[13][31] ) );
  DLH_X1 \bank_register_reg[13][30]  ( .G(n3105), .D(n3234), .Q(
        \bank_register[13][30] ) );
  DLH_X1 \bank_register_reg[13][29]  ( .G(n3103), .D(n3231), .Q(
        \bank_register[13][29] ) );
  DLH_X1 \bank_register_reg[13][28]  ( .G(n3103), .D(n3228), .Q(
        \bank_register[13][28] ) );
  DLH_X1 \bank_register_reg[13][27]  ( .G(n3103), .D(n3225), .Q(
        \bank_register[13][27] ) );
  DLH_X1 \bank_register_reg[13][26]  ( .G(n3103), .D(n3222), .Q(
        \bank_register[13][26] ) );
  DLH_X1 \bank_register_reg[13][25]  ( .G(n3103), .D(n3219), .Q(
        \bank_register[13][25] ) );
  DLH_X1 \bank_register_reg[13][24]  ( .G(n3103), .D(n3216), .Q(
        \bank_register[13][24] ) );
  DLH_X1 \bank_register_reg[13][23]  ( .G(n3103), .D(n3213), .Q(
        \bank_register[13][23] ) );
  DLH_X1 \bank_register_reg[13][22]  ( .G(n3103), .D(n3210), .Q(
        \bank_register[13][22] ) );
  DLH_X1 \bank_register_reg[13][21]  ( .G(n3103), .D(n3207), .Q(
        \bank_register[13][21] ) );
  DLH_X1 \bank_register_reg[13][20]  ( .G(n3103), .D(n3204), .Q(
        \bank_register[13][20] ) );
  DLH_X1 \bank_register_reg[13][19]  ( .G(n3104), .D(n3201), .Q(
        \bank_register[13][19] ) );
  DLH_X1 \bank_register_reg[13][18]  ( .G(n3104), .D(n3198), .Q(
        \bank_register[13][18] ) );
  DLH_X1 \bank_register_reg[13][17]  ( .G(n3105), .D(n3195), .Q(
        \bank_register[13][17] ) );
  DLH_X1 \bank_register_reg[13][16]  ( .G(n3105), .D(n3192), .Q(
        \bank_register[13][16] ) );
  DLH_X1 \bank_register_reg[13][15]  ( .G(n3105), .D(n3189), .Q(
        \bank_register[13][15] ) );
  DLH_X1 \bank_register_reg[13][14]  ( .G(n3105), .D(n3186), .Q(
        \bank_register[13][14] ) );
  DLH_X1 \bank_register_reg[13][13]  ( .G(n3105), .D(n3183), .Q(
        \bank_register[13][13] ) );
  DLH_X1 \bank_register_reg[13][12]  ( .G(n3105), .D(n3180), .Q(
        \bank_register[13][12] ) );
  DLH_X1 \bank_register_reg[13][11]  ( .G(n3105), .D(n3177), .Q(
        \bank_register[13][11] ) );
  DLH_X1 \bank_register_reg[13][10]  ( .G(n3105), .D(n3174), .Q(
        \bank_register[13][10] ) );
  DLH_X1 \bank_register_reg[13][9]  ( .G(n3104), .D(n3171), .Q(
        \bank_register[13][9] ) );
  DLH_X1 \bank_register_reg[13][8]  ( .G(n3104), .D(n3168), .Q(
        \bank_register[13][8] ) );
  DLH_X1 \bank_register_reg[13][7]  ( .G(n3104), .D(n3165), .Q(
        \bank_register[13][7] ) );
  DLH_X1 \bank_register_reg[13][6]  ( .G(n3104), .D(n3162), .Q(
        \bank_register[13][6] ) );
  DLH_X1 \bank_register_reg[13][5]  ( .G(n3104), .D(n3159), .Q(
        \bank_register[13][5] ) );
  DLH_X1 \bank_register_reg[13][4]  ( .G(n3104), .D(n3156), .Q(
        \bank_register[13][4] ) );
  DLH_X1 \bank_register_reg[13][3]  ( .G(n3104), .D(n3153), .Q(
        \bank_register[13][3] ) );
  DLH_X1 \bank_register_reg[13][2]  ( .G(n3104), .D(n3150), .Q(
        \bank_register[13][2] ) );
  DLH_X1 \bank_register_reg[13][1]  ( .G(n3104), .D(n3147), .Q(
        \bank_register[13][1] ) );
  DLH_X1 \bank_register_reg[13][0]  ( .G(n3103), .D(n3144), .Q(
        \bank_register[13][0] ) );
  DLH_X1 \bank_register_reg[14][31]  ( .G(n3102), .D(n3237), .Q(
        \bank_register[14][31] ) );
  DLH_X1 \bank_register_reg[14][30]  ( .G(n3102), .D(n3234), .Q(
        \bank_register[14][30] ) );
  DLH_X1 \bank_register_reg[14][29]  ( .G(n3100), .D(n3231), .Q(
        \bank_register[14][29] ) );
  DLH_X1 \bank_register_reg[14][28]  ( .G(n3100), .D(n3228), .Q(
        \bank_register[14][28] ) );
  DLH_X1 \bank_register_reg[14][27]  ( .G(n3100), .D(n3225), .Q(
        \bank_register[14][27] ) );
  DLH_X1 \bank_register_reg[14][26]  ( .G(n3100), .D(n3222), .Q(
        \bank_register[14][26] ) );
  DLH_X1 \bank_register_reg[14][25]  ( .G(n3100), .D(n3219), .Q(
        \bank_register[14][25] ) );
  DLH_X1 \bank_register_reg[14][24]  ( .G(n3100), .D(n3216), .Q(
        \bank_register[14][24] ) );
  DLH_X1 \bank_register_reg[14][23]  ( .G(n3100), .D(n3213), .Q(
        \bank_register[14][23] ) );
  DLH_X1 \bank_register_reg[14][22]  ( .G(n3100), .D(n3210), .Q(
        \bank_register[14][22] ) );
  DLH_X1 \bank_register_reg[14][21]  ( .G(n3100), .D(n3207), .Q(
        \bank_register[14][21] ) );
  DLH_X1 \bank_register_reg[14][20]  ( .G(n3100), .D(n3204), .Q(
        \bank_register[14][20] ) );
  DLH_X1 \bank_register_reg[14][19]  ( .G(n3101), .D(n3201), .Q(
        \bank_register[14][19] ) );
  DLH_X1 \bank_register_reg[14][18]  ( .G(n3101), .D(n3198), .Q(
        \bank_register[14][18] ) );
  DLH_X1 \bank_register_reg[14][17]  ( .G(n3102), .D(n3195), .Q(
        \bank_register[14][17] ) );
  DLH_X1 \bank_register_reg[14][16]  ( .G(n3102), .D(n3192), .Q(
        \bank_register[14][16] ) );
  DLH_X1 \bank_register_reg[14][15]  ( .G(n3102), .D(n3189), .Q(
        \bank_register[14][15] ) );
  DLH_X1 \bank_register_reg[14][14]  ( .G(n3102), .D(n3186), .Q(
        \bank_register[14][14] ) );
  DLH_X1 \bank_register_reg[14][13]  ( .G(n3102), .D(n3183), .Q(
        \bank_register[14][13] ) );
  DLH_X1 \bank_register_reg[14][12]  ( .G(n3102), .D(n3180), .Q(
        \bank_register[14][12] ) );
  DLH_X1 \bank_register_reg[14][11]  ( .G(n3102), .D(n3177), .Q(
        \bank_register[14][11] ) );
  DLH_X1 \bank_register_reg[14][10]  ( .G(n3102), .D(n3174), .Q(
        \bank_register[14][10] ) );
  DLH_X1 \bank_register_reg[14][9]  ( .G(n3101), .D(n3171), .Q(
        \bank_register[14][9] ) );
  DLH_X1 \bank_register_reg[14][8]  ( .G(n3101), .D(n3168), .Q(
        \bank_register[14][8] ) );
  DLH_X1 \bank_register_reg[14][7]  ( .G(n3101), .D(n3165), .Q(
        \bank_register[14][7] ) );
  DLH_X1 \bank_register_reg[14][6]  ( .G(n3101), .D(n3162), .Q(
        \bank_register[14][6] ) );
  DLH_X1 \bank_register_reg[14][5]  ( .G(n3101), .D(n3159), .Q(
        \bank_register[14][5] ) );
  DLH_X1 \bank_register_reg[14][4]  ( .G(n3101), .D(n3156), .Q(
        \bank_register[14][4] ) );
  DLH_X1 \bank_register_reg[14][3]  ( .G(n3101), .D(n3153), .Q(
        \bank_register[14][3] ) );
  DLH_X1 \bank_register_reg[14][2]  ( .G(n3101), .D(n3150), .Q(
        \bank_register[14][2] ) );
  DLH_X1 \bank_register_reg[14][1]  ( .G(n3101), .D(n3147), .Q(
        \bank_register[14][1] ) );
  DLH_X1 \bank_register_reg[14][0]  ( .G(n3100), .D(n3144), .Q(
        \bank_register[14][0] ) );
  DLH_X1 \bank_register_reg[15][31]  ( .G(n3099), .D(n3237), .Q(
        \bank_register[15][31] ) );
  DLH_X1 \bank_register_reg[15][30]  ( .G(n3099), .D(n3234), .Q(
        \bank_register[15][30] ) );
  DLH_X1 \bank_register_reg[15][29]  ( .G(n3097), .D(n3231), .Q(
        \bank_register[15][29] ) );
  DLH_X1 \bank_register_reg[15][28]  ( .G(n3097), .D(n3228), .Q(
        \bank_register[15][28] ) );
  DLH_X1 \bank_register_reg[15][27]  ( .G(n3097), .D(n3225), .Q(
        \bank_register[15][27] ) );
  DLH_X1 \bank_register_reg[15][26]  ( .G(n3097), .D(n3222), .Q(
        \bank_register[15][26] ) );
  DLH_X1 \bank_register_reg[15][25]  ( .G(n3097), .D(n3219), .Q(
        \bank_register[15][25] ) );
  DLH_X1 \bank_register_reg[15][24]  ( .G(n3097), .D(n3216), .Q(
        \bank_register[15][24] ) );
  DLH_X1 \bank_register_reg[15][23]  ( .G(n3097), .D(n3213), .Q(
        \bank_register[15][23] ) );
  DLH_X1 \bank_register_reg[15][22]  ( .G(n3097), .D(n3210), .Q(
        \bank_register[15][22] ) );
  DLH_X1 \bank_register_reg[15][21]  ( .G(n3097), .D(n3207), .Q(
        \bank_register[15][21] ) );
  DLH_X1 \bank_register_reg[15][20]  ( .G(n3097), .D(n3204), .Q(
        \bank_register[15][20] ) );
  DLH_X1 \bank_register_reg[15][19]  ( .G(n3098), .D(n3201), .Q(
        \bank_register[15][19] ) );
  DLH_X1 \bank_register_reg[15][18]  ( .G(n3098), .D(n3198), .Q(
        \bank_register[15][18] ) );
  DLH_X1 \bank_register_reg[15][17]  ( .G(n3099), .D(n3195), .Q(
        \bank_register[15][17] ) );
  DLH_X1 \bank_register_reg[15][16]  ( .G(n3099), .D(n3192), .Q(
        \bank_register[15][16] ) );
  DLH_X1 \bank_register_reg[15][15]  ( .G(n3099), .D(n3189), .Q(
        \bank_register[15][15] ) );
  DLH_X1 \bank_register_reg[15][14]  ( .G(n3099), .D(n3186), .Q(
        \bank_register[15][14] ) );
  DLH_X1 \bank_register_reg[15][13]  ( .G(n3099), .D(n3183), .Q(
        \bank_register[15][13] ) );
  DLH_X1 \bank_register_reg[15][12]  ( .G(n3099), .D(n3180), .Q(
        \bank_register[15][12] ) );
  DLH_X1 \bank_register_reg[15][11]  ( .G(n3099), .D(n3177), .Q(
        \bank_register[15][11] ) );
  DLH_X1 \bank_register_reg[15][10]  ( .G(n3099), .D(n3174), .Q(
        \bank_register[15][10] ) );
  DLH_X1 \bank_register_reg[15][9]  ( .G(n3098), .D(n3171), .Q(
        \bank_register[15][9] ) );
  DLH_X1 \bank_register_reg[15][8]  ( .G(n3098), .D(n3168), .Q(
        \bank_register[15][8] ) );
  DLH_X1 \bank_register_reg[15][7]  ( .G(n3098), .D(n3165), .Q(
        \bank_register[15][7] ) );
  DLH_X1 \bank_register_reg[15][6]  ( .G(n3098), .D(n3162), .Q(
        \bank_register[15][6] ) );
  DLH_X1 \bank_register_reg[15][5]  ( .G(n3098), .D(n3159), .Q(
        \bank_register[15][5] ) );
  DLH_X1 \bank_register_reg[15][4]  ( .G(n3098), .D(n3156), .Q(
        \bank_register[15][4] ) );
  DLH_X1 \bank_register_reg[15][3]  ( .G(n3098), .D(n3153), .Q(
        \bank_register[15][3] ) );
  DLH_X1 \bank_register_reg[15][2]  ( .G(n3098), .D(n3150), .Q(
        \bank_register[15][2] ) );
  DLH_X1 \bank_register_reg[15][1]  ( .G(n3098), .D(n3147), .Q(
        \bank_register[15][1] ) );
  DLH_X1 \bank_register_reg[15][0]  ( .G(n3097), .D(n3144), .Q(
        \bank_register[15][0] ) );
  DLH_X1 \bank_register_reg[16][31]  ( .G(n3096), .D(n3237), .Q(
        \bank_register[16][31] ) );
  DLH_X1 \bank_register_reg[16][30]  ( .G(n3096), .D(n3234), .Q(
        \bank_register[16][30] ) );
  DLH_X1 \bank_register_reg[16][29]  ( .G(n3094), .D(n3231), .Q(
        \bank_register[16][29] ) );
  DLH_X1 \bank_register_reg[16][28]  ( .G(n3094), .D(n3228), .Q(
        \bank_register[16][28] ) );
  DLH_X1 \bank_register_reg[16][27]  ( .G(n3094), .D(n3225), .Q(
        \bank_register[16][27] ) );
  DLH_X1 \bank_register_reg[16][26]  ( .G(n3094), .D(n3222), .Q(
        \bank_register[16][26] ) );
  DLH_X1 \bank_register_reg[16][25]  ( .G(n3094), .D(n3219), .Q(
        \bank_register[16][25] ) );
  DLH_X1 \bank_register_reg[16][24]  ( .G(n3094), .D(n3216), .Q(
        \bank_register[16][24] ) );
  DLH_X1 \bank_register_reg[16][23]  ( .G(n3094), .D(n3213), .Q(
        \bank_register[16][23] ) );
  DLH_X1 \bank_register_reg[16][22]  ( .G(n3094), .D(n3210), .Q(
        \bank_register[16][22] ) );
  DLH_X1 \bank_register_reg[16][21]  ( .G(n3094), .D(n3207), .Q(
        \bank_register[16][21] ) );
  DLH_X1 \bank_register_reg[16][20]  ( .G(n3094), .D(n3204), .Q(
        \bank_register[16][20] ) );
  DLH_X1 \bank_register_reg[16][19]  ( .G(n3095), .D(n3201), .Q(
        \bank_register[16][19] ) );
  DLH_X1 \bank_register_reg[16][18]  ( .G(n3095), .D(n3198), .Q(
        \bank_register[16][18] ) );
  DLH_X1 \bank_register_reg[16][17]  ( .G(n3096), .D(n3195), .Q(
        \bank_register[16][17] ) );
  DLH_X1 \bank_register_reg[16][16]  ( .G(n3096), .D(n3192), .Q(
        \bank_register[16][16] ) );
  DLH_X1 \bank_register_reg[16][15]  ( .G(n3096), .D(n3189), .Q(
        \bank_register[16][15] ) );
  DLH_X1 \bank_register_reg[16][14]  ( .G(n3096), .D(n3186), .Q(
        \bank_register[16][14] ) );
  DLH_X1 \bank_register_reg[16][13]  ( .G(n3096), .D(n3183), .Q(
        \bank_register[16][13] ) );
  DLH_X1 \bank_register_reg[16][12]  ( .G(n3096), .D(n3180), .Q(
        \bank_register[16][12] ) );
  DLH_X1 \bank_register_reg[16][11]  ( .G(n3096), .D(n3177), .Q(
        \bank_register[16][11] ) );
  DLH_X1 \bank_register_reg[16][10]  ( .G(n3096), .D(n3174), .Q(
        \bank_register[16][10] ) );
  DLH_X1 \bank_register_reg[16][9]  ( .G(n3095), .D(n3171), .Q(
        \bank_register[16][9] ) );
  DLH_X1 \bank_register_reg[16][8]  ( .G(n3095), .D(n3168), .Q(
        \bank_register[16][8] ) );
  DLH_X1 \bank_register_reg[16][7]  ( .G(n3095), .D(n3165), .Q(
        \bank_register[16][7] ) );
  DLH_X1 \bank_register_reg[16][6]  ( .G(n3095), .D(n3162), .Q(
        \bank_register[16][6] ) );
  DLH_X1 \bank_register_reg[16][5]  ( .G(n3095), .D(n3159), .Q(
        \bank_register[16][5] ) );
  DLH_X1 \bank_register_reg[16][4]  ( .G(n3095), .D(n3156), .Q(
        \bank_register[16][4] ) );
  DLH_X1 \bank_register_reg[16][3]  ( .G(n3095), .D(n3153), .Q(
        \bank_register[16][3] ) );
  DLH_X1 \bank_register_reg[16][2]  ( .G(n3095), .D(n3150), .Q(
        \bank_register[16][2] ) );
  DLH_X1 \bank_register_reg[16][1]  ( .G(n3095), .D(n3147), .Q(
        \bank_register[16][1] ) );
  DLH_X1 \bank_register_reg[16][0]  ( .G(n3094), .D(n3144), .Q(
        \bank_register[16][0] ) );
  DLH_X1 \bank_register_reg[17][31]  ( .G(n3093), .D(n3237), .Q(
        \bank_register[17][31] ) );
  DLH_X1 \bank_register_reg[17][30]  ( .G(n3093), .D(n3234), .Q(
        \bank_register[17][30] ) );
  DLH_X1 \bank_register_reg[17][29]  ( .G(n3091), .D(n3231), .Q(
        \bank_register[17][29] ) );
  DLH_X1 \bank_register_reg[17][28]  ( .G(n3091), .D(n3228), .Q(
        \bank_register[17][28] ) );
  DLH_X1 \bank_register_reg[17][27]  ( .G(n3091), .D(n3225), .Q(
        \bank_register[17][27] ) );
  DLH_X1 \bank_register_reg[17][26]  ( .G(n3091), .D(n3222), .Q(
        \bank_register[17][26] ) );
  DLH_X1 \bank_register_reg[17][25]  ( .G(n3091), .D(n3219), .Q(
        \bank_register[17][25] ) );
  DLH_X1 \bank_register_reg[17][24]  ( .G(n3091), .D(n3216), .Q(
        \bank_register[17][24] ) );
  DLH_X1 \bank_register_reg[17][23]  ( .G(n3091), .D(n3213), .Q(
        \bank_register[17][23] ) );
  DLH_X1 \bank_register_reg[17][22]  ( .G(n3091), .D(n3210), .Q(
        \bank_register[17][22] ) );
  DLH_X1 \bank_register_reg[17][21]  ( .G(n3091), .D(n3207), .Q(
        \bank_register[17][21] ) );
  DLH_X1 \bank_register_reg[17][20]  ( .G(n3091), .D(n3204), .Q(
        \bank_register[17][20] ) );
  DLH_X1 \bank_register_reg[17][19]  ( .G(n3092), .D(n3201), .Q(
        \bank_register[17][19] ) );
  DLH_X1 \bank_register_reg[17][18]  ( .G(n3092), .D(n3198), .Q(
        \bank_register[17][18] ) );
  DLH_X1 \bank_register_reg[17][17]  ( .G(n3093), .D(n3195), .Q(
        \bank_register[17][17] ) );
  DLH_X1 \bank_register_reg[17][16]  ( .G(n3093), .D(n3192), .Q(
        \bank_register[17][16] ) );
  DLH_X1 \bank_register_reg[17][15]  ( .G(n3093), .D(n3189), .Q(
        \bank_register[17][15] ) );
  DLH_X1 \bank_register_reg[17][14]  ( .G(n3093), .D(n3186), .Q(
        \bank_register[17][14] ) );
  DLH_X1 \bank_register_reg[17][13]  ( .G(n3093), .D(n3183), .Q(
        \bank_register[17][13] ) );
  DLH_X1 \bank_register_reg[17][12]  ( .G(n3093), .D(n3180), .Q(
        \bank_register[17][12] ) );
  DLH_X1 \bank_register_reg[17][11]  ( .G(n3093), .D(n3177), .Q(
        \bank_register[17][11] ) );
  DLH_X1 \bank_register_reg[17][10]  ( .G(n3093), .D(n3174), .Q(
        \bank_register[17][10] ) );
  DLH_X1 \bank_register_reg[17][9]  ( .G(n3092), .D(n3171), .Q(
        \bank_register[17][9] ) );
  DLH_X1 \bank_register_reg[17][8]  ( .G(n3092), .D(n3168), .Q(
        \bank_register[17][8] ) );
  DLH_X1 \bank_register_reg[17][7]  ( .G(n3092), .D(n3165), .Q(
        \bank_register[17][7] ) );
  DLH_X1 \bank_register_reg[17][6]  ( .G(n3092), .D(n3162), .Q(
        \bank_register[17][6] ) );
  DLH_X1 \bank_register_reg[17][5]  ( .G(n3092), .D(n3159), .Q(
        \bank_register[17][5] ) );
  DLH_X1 \bank_register_reg[17][4]  ( .G(n3092), .D(n3156), .Q(
        \bank_register[17][4] ) );
  DLH_X1 \bank_register_reg[17][3]  ( .G(n3092), .D(n3153), .Q(
        \bank_register[17][3] ) );
  DLH_X1 \bank_register_reg[17][2]  ( .G(n3092), .D(n3150), .Q(
        \bank_register[17][2] ) );
  DLH_X1 \bank_register_reg[17][1]  ( .G(n3092), .D(n3147), .Q(
        \bank_register[17][1] ) );
  DLH_X1 \bank_register_reg[17][0]  ( .G(n3091), .D(n3144), .Q(
        \bank_register[17][0] ) );
  DLH_X1 \bank_register_reg[18][31]  ( .G(n3090), .D(n3237), .Q(
        \bank_register[18][31] ) );
  DLH_X1 \bank_register_reg[18][30]  ( .G(n3090), .D(n3234), .Q(
        \bank_register[18][30] ) );
  DLH_X1 \bank_register_reg[18][29]  ( .G(n3088), .D(n3231), .Q(
        \bank_register[18][29] ) );
  DLH_X1 \bank_register_reg[18][28]  ( .G(n3088), .D(n3228), .Q(
        \bank_register[18][28] ) );
  DLH_X1 \bank_register_reg[18][27]  ( .G(n3088), .D(n3225), .Q(
        \bank_register[18][27] ) );
  DLH_X1 \bank_register_reg[18][26]  ( .G(n3088), .D(n3222), .Q(
        \bank_register[18][26] ) );
  DLH_X1 \bank_register_reg[18][25]  ( .G(n3088), .D(n3219), .Q(
        \bank_register[18][25] ) );
  DLH_X1 \bank_register_reg[18][24]  ( .G(n3088), .D(n3216), .Q(
        \bank_register[18][24] ) );
  DLH_X1 \bank_register_reg[18][23]  ( .G(n3088), .D(n3213), .Q(
        \bank_register[18][23] ) );
  DLH_X1 \bank_register_reg[18][22]  ( .G(n3088), .D(n3210), .Q(
        \bank_register[18][22] ) );
  DLH_X1 \bank_register_reg[18][21]  ( .G(n3088), .D(n3207), .Q(
        \bank_register[18][21] ) );
  DLH_X1 \bank_register_reg[18][20]  ( .G(n3088), .D(n3204), .Q(
        \bank_register[18][20] ) );
  DLH_X1 \bank_register_reg[18][19]  ( .G(n3089), .D(n3201), .Q(
        \bank_register[18][19] ) );
  DLH_X1 \bank_register_reg[18][18]  ( .G(n3089), .D(n3198), .Q(
        \bank_register[18][18] ) );
  DLH_X1 \bank_register_reg[18][17]  ( .G(n3090), .D(n3195), .Q(
        \bank_register[18][17] ) );
  DLH_X1 \bank_register_reg[18][16]  ( .G(n3090), .D(n3192), .Q(
        \bank_register[18][16] ) );
  DLH_X1 \bank_register_reg[18][15]  ( .G(n3090), .D(n3189), .Q(
        \bank_register[18][15] ) );
  DLH_X1 \bank_register_reg[18][14]  ( .G(n3090), .D(n3186), .Q(
        \bank_register[18][14] ) );
  DLH_X1 \bank_register_reg[18][13]  ( .G(n3090), .D(n3183), .Q(
        \bank_register[18][13] ) );
  DLH_X1 \bank_register_reg[18][12]  ( .G(n3090), .D(n3180), .Q(
        \bank_register[18][12] ) );
  DLH_X1 \bank_register_reg[18][11]  ( .G(n3090), .D(n3177), .Q(
        \bank_register[18][11] ) );
  DLH_X1 \bank_register_reg[18][10]  ( .G(n3090), .D(n3174), .Q(
        \bank_register[18][10] ) );
  DLH_X1 \bank_register_reg[18][9]  ( .G(n3089), .D(n3171), .Q(
        \bank_register[18][9] ) );
  DLH_X1 \bank_register_reg[18][8]  ( .G(n3089), .D(n3168), .Q(
        \bank_register[18][8] ) );
  DLH_X1 \bank_register_reg[18][7]  ( .G(n3089), .D(n3165), .Q(
        \bank_register[18][7] ) );
  DLH_X1 \bank_register_reg[18][6]  ( .G(n3089), .D(n3162), .Q(
        \bank_register[18][6] ) );
  DLH_X1 \bank_register_reg[18][5]  ( .G(n3089), .D(n3159), .Q(
        \bank_register[18][5] ) );
  DLH_X1 \bank_register_reg[18][4]  ( .G(n3089), .D(n3156), .Q(
        \bank_register[18][4] ) );
  DLH_X1 \bank_register_reg[18][3]  ( .G(n3089), .D(n3153), .Q(
        \bank_register[18][3] ) );
  DLH_X1 \bank_register_reg[18][2]  ( .G(n3089), .D(n3150), .Q(
        \bank_register[18][2] ) );
  DLH_X1 \bank_register_reg[18][1]  ( .G(n3089), .D(n3147), .Q(
        \bank_register[18][1] ) );
  DLH_X1 \bank_register_reg[18][0]  ( .G(n3088), .D(n3144), .Q(
        \bank_register[18][0] ) );
  DLH_X1 \bank_register_reg[19][31]  ( .G(n3087), .D(n3237), .Q(
        \bank_register[19][31] ) );
  DLH_X1 \bank_register_reg[19][30]  ( .G(n3087), .D(n3234), .Q(
        \bank_register[19][30] ) );
  DLH_X1 \bank_register_reg[19][29]  ( .G(n3085), .D(n3231), .Q(
        \bank_register[19][29] ) );
  DLH_X1 \bank_register_reg[19][28]  ( .G(n3085), .D(n3228), .Q(
        \bank_register[19][28] ) );
  DLH_X1 \bank_register_reg[19][27]  ( .G(n3085), .D(n3225), .Q(
        \bank_register[19][27] ) );
  DLH_X1 \bank_register_reg[19][26]  ( .G(n3085), .D(n3222), .Q(
        \bank_register[19][26] ) );
  DLH_X1 \bank_register_reg[19][25]  ( .G(n3085), .D(n3219), .Q(
        \bank_register[19][25] ) );
  DLH_X1 \bank_register_reg[19][24]  ( .G(n3085), .D(n3216), .Q(
        \bank_register[19][24] ) );
  DLH_X1 \bank_register_reg[19][23]  ( .G(n3085), .D(n3213), .Q(
        \bank_register[19][23] ) );
  DLH_X1 \bank_register_reg[19][22]  ( .G(n3085), .D(n3210), .Q(
        \bank_register[19][22] ) );
  DLH_X1 \bank_register_reg[19][21]  ( .G(n3085), .D(n3207), .Q(
        \bank_register[19][21] ) );
  DLH_X1 \bank_register_reg[19][20]  ( .G(n3085), .D(n3204), .Q(
        \bank_register[19][20] ) );
  DLH_X1 \bank_register_reg[19][19]  ( .G(n3086), .D(n3201), .Q(
        \bank_register[19][19] ) );
  DLH_X1 \bank_register_reg[19][18]  ( .G(n3086), .D(n3198), .Q(
        \bank_register[19][18] ) );
  DLH_X1 \bank_register_reg[19][17]  ( .G(n3087), .D(n3195), .Q(
        \bank_register[19][17] ) );
  DLH_X1 \bank_register_reg[19][16]  ( .G(n3087), .D(n3192), .Q(
        \bank_register[19][16] ) );
  DLH_X1 \bank_register_reg[19][15]  ( .G(n3087), .D(n3189), .Q(
        \bank_register[19][15] ) );
  DLH_X1 \bank_register_reg[19][14]  ( .G(n3087), .D(n3186), .Q(
        \bank_register[19][14] ) );
  DLH_X1 \bank_register_reg[19][13]  ( .G(n3087), .D(n3183), .Q(
        \bank_register[19][13] ) );
  DLH_X1 \bank_register_reg[19][12]  ( .G(n3087), .D(n3180), .Q(
        \bank_register[19][12] ) );
  DLH_X1 \bank_register_reg[19][11]  ( .G(n3087), .D(n3177), .Q(
        \bank_register[19][11] ) );
  DLH_X1 \bank_register_reg[19][10]  ( .G(n3087), .D(n3174), .Q(
        \bank_register[19][10] ) );
  DLH_X1 \bank_register_reg[19][9]  ( .G(n3086), .D(n3171), .Q(
        \bank_register[19][9] ) );
  DLH_X1 \bank_register_reg[19][8]  ( .G(n3086), .D(n3168), .Q(
        \bank_register[19][8] ) );
  DLH_X1 \bank_register_reg[19][7]  ( .G(n3086), .D(n3165), .Q(
        \bank_register[19][7] ) );
  DLH_X1 \bank_register_reg[19][6]  ( .G(n3086), .D(n3162), .Q(
        \bank_register[19][6] ) );
  DLH_X1 \bank_register_reg[19][5]  ( .G(n3086), .D(n3159), .Q(
        \bank_register[19][5] ) );
  DLH_X1 \bank_register_reg[19][4]  ( .G(n3086), .D(n3156), .Q(
        \bank_register[19][4] ) );
  DLH_X1 \bank_register_reg[19][3]  ( .G(n3086), .D(n3153), .Q(
        \bank_register[19][3] ) );
  DLH_X1 \bank_register_reg[19][2]  ( .G(n3086), .D(n3150), .Q(
        \bank_register[19][2] ) );
  DLH_X1 \bank_register_reg[19][1]  ( .G(n3086), .D(n3147), .Q(
        \bank_register[19][1] ) );
  DLH_X1 \bank_register_reg[19][0]  ( .G(n3085), .D(n3144), .Q(
        \bank_register[19][0] ) );
  DLH_X1 \bank_register_reg[20][31]  ( .G(n3084), .D(n3236), .Q(
        \bank_register[20][31] ) );
  DLH_X1 \bank_register_reg[20][30]  ( .G(n3084), .D(n3233), .Q(
        \bank_register[20][30] ) );
  DLH_X1 \bank_register_reg[20][29]  ( .G(n3082), .D(n3230), .Q(
        \bank_register[20][29] ) );
  DLH_X1 \bank_register_reg[20][28]  ( .G(n3082), .D(n3227), .Q(
        \bank_register[20][28] ) );
  DLH_X1 \bank_register_reg[20][27]  ( .G(n3082), .D(n3224), .Q(
        \bank_register[20][27] ) );
  DLH_X1 \bank_register_reg[20][26]  ( .G(n3082), .D(n3221), .Q(
        \bank_register[20][26] ) );
  DLH_X1 \bank_register_reg[20][25]  ( .G(n3082), .D(n3218), .Q(
        \bank_register[20][25] ) );
  DLH_X1 \bank_register_reg[20][24]  ( .G(n3082), .D(n3215), .Q(
        \bank_register[20][24] ) );
  DLH_X1 \bank_register_reg[20][23]  ( .G(n3082), .D(n3212), .Q(
        \bank_register[20][23] ) );
  DLH_X1 \bank_register_reg[20][22]  ( .G(n3082), .D(n3209), .Q(
        \bank_register[20][22] ) );
  DLH_X1 \bank_register_reg[20][21]  ( .G(n3082), .D(n3206), .Q(
        \bank_register[20][21] ) );
  DLH_X1 \bank_register_reg[20][20]  ( .G(n3082), .D(n3203), .Q(
        \bank_register[20][20] ) );
  DLH_X1 \bank_register_reg[20][19]  ( .G(n3083), .D(n3200), .Q(
        \bank_register[20][19] ) );
  DLH_X1 \bank_register_reg[20][18]  ( .G(n3083), .D(n3197), .Q(
        \bank_register[20][18] ) );
  DLH_X1 \bank_register_reg[20][17]  ( .G(n3084), .D(n3194), .Q(
        \bank_register[20][17] ) );
  DLH_X1 \bank_register_reg[20][16]  ( .G(n3084), .D(n3191), .Q(
        \bank_register[20][16] ) );
  DLH_X1 \bank_register_reg[20][15]  ( .G(n3084), .D(n3188), .Q(
        \bank_register[20][15] ) );
  DLH_X1 \bank_register_reg[20][14]  ( .G(n3084), .D(n3185), .Q(
        \bank_register[20][14] ) );
  DLH_X1 \bank_register_reg[20][13]  ( .G(n3084), .D(n3182), .Q(
        \bank_register[20][13] ) );
  DLH_X1 \bank_register_reg[20][12]  ( .G(n3084), .D(n3179), .Q(
        \bank_register[20][12] ) );
  DLH_X1 \bank_register_reg[20][11]  ( .G(n3084), .D(n3176), .Q(
        \bank_register[20][11] ) );
  DLH_X1 \bank_register_reg[20][10]  ( .G(n3084), .D(n3173), .Q(
        \bank_register[20][10] ) );
  DLH_X1 \bank_register_reg[20][9]  ( .G(n3083), .D(n3170), .Q(
        \bank_register[20][9] ) );
  DLH_X1 \bank_register_reg[20][8]  ( .G(n3083), .D(n3167), .Q(
        \bank_register[20][8] ) );
  DLH_X1 \bank_register_reg[20][7]  ( .G(n3083), .D(n3164), .Q(
        \bank_register[20][7] ) );
  DLH_X1 \bank_register_reg[20][6]  ( .G(n3083), .D(n3161), .Q(
        \bank_register[20][6] ) );
  DLH_X1 \bank_register_reg[20][5]  ( .G(n3083), .D(n3158), .Q(
        \bank_register[20][5] ) );
  DLH_X1 \bank_register_reg[20][4]  ( .G(n3083), .D(n3155), .Q(
        \bank_register[20][4] ) );
  DLH_X1 \bank_register_reg[20][3]  ( .G(n3083), .D(n3152), .Q(
        \bank_register[20][3] ) );
  DLH_X1 \bank_register_reg[20][2]  ( .G(n3083), .D(n3149), .Q(
        \bank_register[20][2] ) );
  DLH_X1 \bank_register_reg[20][1]  ( .G(n3083), .D(n3146), .Q(
        \bank_register[20][1] ) );
  DLH_X1 \bank_register_reg[20][0]  ( .G(n3082), .D(n3143), .Q(
        \bank_register[20][0] ) );
  DLH_X1 \bank_register_reg[21][31]  ( .G(n3081), .D(n3235), .Q(
        \bank_register[21][31] ) );
  DLH_X1 \bank_register_reg[21][30]  ( .G(n3081), .D(n3232), .Q(
        \bank_register[21][30] ) );
  DLH_X1 \bank_register_reg[21][29]  ( .G(n3079), .D(n3229), .Q(
        \bank_register[21][29] ) );
  DLH_X1 \bank_register_reg[21][28]  ( .G(n3079), .D(n3226), .Q(
        \bank_register[21][28] ) );
  DLH_X1 \bank_register_reg[21][27]  ( .G(n3079), .D(n3223), .Q(
        \bank_register[21][27] ) );
  DLH_X1 \bank_register_reg[21][26]  ( .G(n3079), .D(n3220), .Q(
        \bank_register[21][26] ) );
  DLH_X1 \bank_register_reg[21][25]  ( .G(n3079), .D(n3217), .Q(
        \bank_register[21][25] ) );
  DLH_X1 \bank_register_reg[21][24]  ( .G(n3079), .D(n3214), .Q(
        \bank_register[21][24] ) );
  DLH_X1 \bank_register_reg[21][23]  ( .G(n3079), .D(n3211), .Q(
        \bank_register[21][23] ) );
  DLH_X1 \bank_register_reg[21][22]  ( .G(n3079), .D(n3208), .Q(
        \bank_register[21][22] ) );
  DLH_X1 \bank_register_reg[21][21]  ( .G(n3079), .D(n3205), .Q(
        \bank_register[21][21] ) );
  DLH_X1 \bank_register_reg[21][20]  ( .G(n3079), .D(n3202), .Q(
        \bank_register[21][20] ) );
  DLH_X1 \bank_register_reg[21][19]  ( .G(n3080), .D(n3199), .Q(
        \bank_register[21][19] ) );
  DLH_X1 \bank_register_reg[21][18]  ( .G(n3080), .D(n3196), .Q(
        \bank_register[21][18] ) );
  DLH_X1 \bank_register_reg[21][17]  ( .G(n3081), .D(n3193), .Q(
        \bank_register[21][17] ) );
  DLH_X1 \bank_register_reg[21][16]  ( .G(n3081), .D(n3190), .Q(
        \bank_register[21][16] ) );
  DLH_X1 \bank_register_reg[21][15]  ( .G(n3081), .D(n3187), .Q(
        \bank_register[21][15] ) );
  DLH_X1 \bank_register_reg[21][14]  ( .G(n3081), .D(n3184), .Q(
        \bank_register[21][14] ) );
  DLH_X1 \bank_register_reg[21][13]  ( .G(n3081), .D(n3181), .Q(
        \bank_register[21][13] ) );
  DLH_X1 \bank_register_reg[21][12]  ( .G(n3081), .D(n3178), .Q(
        \bank_register[21][12] ) );
  DLH_X1 \bank_register_reg[21][11]  ( .G(n3081), .D(n3175), .Q(
        \bank_register[21][11] ) );
  DLH_X1 \bank_register_reg[21][10]  ( .G(n3081), .D(n3172), .Q(
        \bank_register[21][10] ) );
  DLH_X1 \bank_register_reg[21][9]  ( .G(n3080), .D(n3169), .Q(
        \bank_register[21][9] ) );
  DLH_X1 \bank_register_reg[21][8]  ( .G(n3080), .D(n3166), .Q(
        \bank_register[21][8] ) );
  DLH_X1 \bank_register_reg[21][7]  ( .G(n3080), .D(n3163), .Q(
        \bank_register[21][7] ) );
  DLH_X1 \bank_register_reg[21][6]  ( .G(n3080), .D(n3160), .Q(
        \bank_register[21][6] ) );
  DLH_X1 \bank_register_reg[21][5]  ( .G(n3080), .D(n3157), .Q(
        \bank_register[21][5] ) );
  DLH_X1 \bank_register_reg[21][4]  ( .G(n3080), .D(n3154), .Q(
        \bank_register[21][4] ) );
  DLH_X1 \bank_register_reg[21][3]  ( .G(n3080), .D(n3151), .Q(
        \bank_register[21][3] ) );
  DLH_X1 \bank_register_reg[21][2]  ( .G(n3080), .D(n3148), .Q(
        \bank_register[21][2] ) );
  DLH_X1 \bank_register_reg[21][1]  ( .G(n3080), .D(n3145), .Q(
        \bank_register[21][1] ) );
  DLH_X1 \bank_register_reg[21][0]  ( .G(n3079), .D(n3142), .Q(
        \bank_register[21][0] ) );
  DLH_X1 \bank_register_reg[22][31]  ( .G(n3078), .D(n3235), .Q(
        \bank_register[22][31] ) );
  DLH_X1 \bank_register_reg[22][30]  ( .G(n3078), .D(n3232), .Q(
        \bank_register[22][30] ) );
  DLH_X1 \bank_register_reg[22][29]  ( .G(n3076), .D(n3229), .Q(
        \bank_register[22][29] ) );
  DLH_X1 \bank_register_reg[22][28]  ( .G(n3076), .D(n3226), .Q(
        \bank_register[22][28] ) );
  DLH_X1 \bank_register_reg[22][27]  ( .G(n3076), .D(n3223), .Q(
        \bank_register[22][27] ) );
  DLH_X1 \bank_register_reg[22][26]  ( .G(n3076), .D(n3220), .Q(
        \bank_register[22][26] ) );
  DLH_X1 \bank_register_reg[22][25]  ( .G(n3076), .D(n3217), .Q(
        \bank_register[22][25] ) );
  DLH_X1 \bank_register_reg[22][24]  ( .G(n3076), .D(n3214), .Q(
        \bank_register[22][24] ) );
  DLH_X1 \bank_register_reg[22][23]  ( .G(n3076), .D(n3211), .Q(
        \bank_register[22][23] ) );
  DLH_X1 \bank_register_reg[22][22]  ( .G(n3076), .D(n3208), .Q(
        \bank_register[22][22] ) );
  DLH_X1 \bank_register_reg[22][21]  ( .G(n3076), .D(n3205), .Q(
        \bank_register[22][21] ) );
  DLH_X1 \bank_register_reg[22][20]  ( .G(n3076), .D(n3202), .Q(
        \bank_register[22][20] ) );
  DLH_X1 \bank_register_reg[22][19]  ( .G(n3077), .D(n3199), .Q(
        \bank_register[22][19] ) );
  DLH_X1 \bank_register_reg[22][18]  ( .G(n3077), .D(n3196), .Q(
        \bank_register[22][18] ) );
  DLH_X1 \bank_register_reg[22][17]  ( .G(n3078), .D(n3193), .Q(
        \bank_register[22][17] ) );
  DLH_X1 \bank_register_reg[22][16]  ( .G(n3078), .D(n3190), .Q(
        \bank_register[22][16] ) );
  DLH_X1 \bank_register_reg[22][15]  ( .G(n3078), .D(n3187), .Q(
        \bank_register[22][15] ) );
  DLH_X1 \bank_register_reg[22][14]  ( .G(n3078), .D(n3184), .Q(
        \bank_register[22][14] ) );
  DLH_X1 \bank_register_reg[22][13]  ( .G(n3078), .D(n3181), .Q(
        \bank_register[22][13] ) );
  DLH_X1 \bank_register_reg[22][12]  ( .G(n3078), .D(n3178), .Q(
        \bank_register[22][12] ) );
  DLH_X1 \bank_register_reg[22][11]  ( .G(n3078), .D(n3175), .Q(
        \bank_register[22][11] ) );
  DLH_X1 \bank_register_reg[22][10]  ( .G(n3078), .D(n3172), .Q(
        \bank_register[22][10] ) );
  DLH_X1 \bank_register_reg[22][9]  ( .G(n3077), .D(n3169), .Q(
        \bank_register[22][9] ) );
  DLH_X1 \bank_register_reg[22][8]  ( .G(n3077), .D(n3166), .Q(
        \bank_register[22][8] ) );
  DLH_X1 \bank_register_reg[22][7]  ( .G(n3077), .D(n3163), .Q(
        \bank_register[22][7] ) );
  DLH_X1 \bank_register_reg[22][6]  ( .G(n3077), .D(n3160), .Q(
        \bank_register[22][6] ) );
  DLH_X1 \bank_register_reg[22][5]  ( .G(n3077), .D(n3157), .Q(
        \bank_register[22][5] ) );
  DLH_X1 \bank_register_reg[22][4]  ( .G(n3077), .D(n3154), .Q(
        \bank_register[22][4] ) );
  DLH_X1 \bank_register_reg[22][3]  ( .G(n3077), .D(n3151), .Q(
        \bank_register[22][3] ) );
  DLH_X1 \bank_register_reg[22][2]  ( .G(n3077), .D(n3148), .Q(
        \bank_register[22][2] ) );
  DLH_X1 \bank_register_reg[22][1]  ( .G(n3077), .D(n3145), .Q(
        \bank_register[22][1] ) );
  DLH_X1 \bank_register_reg[22][0]  ( .G(n3076), .D(n3142), .Q(
        \bank_register[22][0] ) );
  DLH_X1 \bank_register_reg[23][31]  ( .G(n3075), .D(n3235), .Q(
        \bank_register[23][31] ) );
  DLH_X1 \bank_register_reg[23][30]  ( .G(n3075), .D(n3232), .Q(
        \bank_register[23][30] ) );
  DLH_X1 \bank_register_reg[23][29]  ( .G(n3073), .D(n3229), .Q(
        \bank_register[23][29] ) );
  DLH_X1 \bank_register_reg[23][28]  ( .G(n3073), .D(n3226), .Q(
        \bank_register[23][28] ) );
  DLH_X1 \bank_register_reg[23][27]  ( .G(n3073), .D(n3223), .Q(
        \bank_register[23][27] ) );
  DLH_X1 \bank_register_reg[23][26]  ( .G(n3073), .D(n3220), .Q(
        \bank_register[23][26] ) );
  DLH_X1 \bank_register_reg[23][25]  ( .G(n3073), .D(n3217), .Q(
        \bank_register[23][25] ) );
  DLH_X1 \bank_register_reg[23][24]  ( .G(n3073), .D(n3214), .Q(
        \bank_register[23][24] ) );
  DLH_X1 \bank_register_reg[23][23]  ( .G(n3073), .D(n3211), .Q(
        \bank_register[23][23] ) );
  DLH_X1 \bank_register_reg[23][22]  ( .G(n3073), .D(n3208), .Q(
        \bank_register[23][22] ) );
  DLH_X1 \bank_register_reg[23][21]  ( .G(n3073), .D(n3205), .Q(
        \bank_register[23][21] ) );
  DLH_X1 \bank_register_reg[23][20]  ( .G(n3073), .D(n3202), .Q(
        \bank_register[23][20] ) );
  DLH_X1 \bank_register_reg[23][19]  ( .G(n3074), .D(n3199), .Q(
        \bank_register[23][19] ) );
  DLH_X1 \bank_register_reg[23][18]  ( .G(n3074), .D(n3196), .Q(
        \bank_register[23][18] ) );
  DLH_X1 \bank_register_reg[23][17]  ( .G(n3075), .D(n3193), .Q(
        \bank_register[23][17] ) );
  DLH_X1 \bank_register_reg[23][16]  ( .G(n3075), .D(n3190), .Q(
        \bank_register[23][16] ) );
  DLH_X1 \bank_register_reg[23][15]  ( .G(n3075), .D(n3187), .Q(
        \bank_register[23][15] ) );
  DLH_X1 \bank_register_reg[23][14]  ( .G(n3075), .D(n3184), .Q(
        \bank_register[23][14] ) );
  DLH_X1 \bank_register_reg[23][13]  ( .G(n3075), .D(n3181), .Q(
        \bank_register[23][13] ) );
  DLH_X1 \bank_register_reg[23][12]  ( .G(n3075), .D(n3178), .Q(
        \bank_register[23][12] ) );
  DLH_X1 \bank_register_reg[23][11]  ( .G(n3075), .D(n3175), .Q(
        \bank_register[23][11] ) );
  DLH_X1 \bank_register_reg[23][10]  ( .G(n3075), .D(n3172), .Q(
        \bank_register[23][10] ) );
  DLH_X1 \bank_register_reg[23][9]  ( .G(n3074), .D(n3169), .Q(
        \bank_register[23][9] ) );
  DLH_X1 \bank_register_reg[23][8]  ( .G(n3074), .D(n3166), .Q(
        \bank_register[23][8] ) );
  DLH_X1 \bank_register_reg[23][7]  ( .G(n3074), .D(n3163), .Q(
        \bank_register[23][7] ) );
  DLH_X1 \bank_register_reg[23][6]  ( .G(n3074), .D(n3160), .Q(
        \bank_register[23][6] ) );
  DLH_X1 \bank_register_reg[23][5]  ( .G(n3074), .D(n3157), .Q(
        \bank_register[23][5] ) );
  DLH_X1 \bank_register_reg[23][4]  ( .G(n3074), .D(n3154), .Q(
        \bank_register[23][4] ) );
  DLH_X1 \bank_register_reg[23][3]  ( .G(n3074), .D(n3151), .Q(
        \bank_register[23][3] ) );
  DLH_X1 \bank_register_reg[23][2]  ( .G(n3074), .D(n3148), .Q(
        \bank_register[23][2] ) );
  DLH_X1 \bank_register_reg[23][1]  ( .G(n3074), .D(n3145), .Q(
        \bank_register[23][1] ) );
  DLH_X1 \bank_register_reg[23][0]  ( .G(n3073), .D(n3142), .Q(
        \bank_register[23][0] ) );
  DLH_X1 \bank_register_reg[24][31]  ( .G(n3072), .D(n3235), .Q(
        \bank_register[24][31] ) );
  DLH_X1 \bank_register_reg[24][30]  ( .G(n3072), .D(n3232), .Q(
        \bank_register[24][30] ) );
  DLH_X1 \bank_register_reg[24][29]  ( .G(n3070), .D(n3229), .Q(
        \bank_register[24][29] ) );
  DLH_X1 \bank_register_reg[24][28]  ( .G(n3070), .D(n3226), .Q(
        \bank_register[24][28] ) );
  DLH_X1 \bank_register_reg[24][27]  ( .G(n3070), .D(n3223), .Q(
        \bank_register[24][27] ) );
  DLH_X1 \bank_register_reg[24][26]  ( .G(n3070), .D(n3220), .Q(
        \bank_register[24][26] ) );
  DLH_X1 \bank_register_reg[24][25]  ( .G(n3070), .D(n3217), .Q(
        \bank_register[24][25] ) );
  DLH_X1 \bank_register_reg[24][24]  ( .G(n3070), .D(n3214), .Q(
        \bank_register[24][24] ) );
  DLH_X1 \bank_register_reg[24][23]  ( .G(n3070), .D(n3211), .Q(
        \bank_register[24][23] ) );
  DLH_X1 \bank_register_reg[24][22]  ( .G(n3070), .D(n3208), .Q(
        \bank_register[24][22] ) );
  DLH_X1 \bank_register_reg[24][21]  ( .G(n3070), .D(n3205), .Q(
        \bank_register[24][21] ) );
  DLH_X1 \bank_register_reg[24][20]  ( .G(n3070), .D(n3202), .Q(
        \bank_register[24][20] ) );
  DLH_X1 \bank_register_reg[24][19]  ( .G(n3071), .D(n3199), .Q(
        \bank_register[24][19] ) );
  DLH_X1 \bank_register_reg[24][18]  ( .G(n3071), .D(n3196), .Q(
        \bank_register[24][18] ) );
  DLH_X1 \bank_register_reg[24][17]  ( .G(n3072), .D(n3193), .Q(
        \bank_register[24][17] ) );
  DLH_X1 \bank_register_reg[24][16]  ( .G(n3072), .D(n3190), .Q(
        \bank_register[24][16] ) );
  DLH_X1 \bank_register_reg[24][15]  ( .G(n3072), .D(n3187), .Q(
        \bank_register[24][15] ) );
  DLH_X1 \bank_register_reg[24][14]  ( .G(n3072), .D(n3184), .Q(
        \bank_register[24][14] ) );
  DLH_X1 \bank_register_reg[24][13]  ( .G(n3072), .D(n3181), .Q(
        \bank_register[24][13] ) );
  DLH_X1 \bank_register_reg[24][12]  ( .G(n3072), .D(n3178), .Q(
        \bank_register[24][12] ) );
  DLH_X1 \bank_register_reg[24][11]  ( .G(n3072), .D(n3175), .Q(
        \bank_register[24][11] ) );
  DLH_X1 \bank_register_reg[24][10]  ( .G(n3072), .D(n3172), .Q(
        \bank_register[24][10] ) );
  DLH_X1 \bank_register_reg[24][9]  ( .G(n3071), .D(n3169), .Q(
        \bank_register[24][9] ) );
  DLH_X1 \bank_register_reg[24][8]  ( .G(n3071), .D(n3166), .Q(
        \bank_register[24][8] ) );
  DLH_X1 \bank_register_reg[24][7]  ( .G(n3071), .D(n3163), .Q(
        \bank_register[24][7] ) );
  DLH_X1 \bank_register_reg[24][6]  ( .G(n3071), .D(n3160), .Q(
        \bank_register[24][6] ) );
  DLH_X1 \bank_register_reg[24][5]  ( .G(n3071), .D(n3157), .Q(
        \bank_register[24][5] ) );
  DLH_X1 \bank_register_reg[24][4]  ( .G(n3071), .D(n3154), .Q(
        \bank_register[24][4] ) );
  DLH_X1 \bank_register_reg[24][3]  ( .G(n3071), .D(n3151), .Q(
        \bank_register[24][3] ) );
  DLH_X1 \bank_register_reg[24][2]  ( .G(n3071), .D(n3148), .Q(
        \bank_register[24][2] ) );
  DLH_X1 \bank_register_reg[24][1]  ( .G(n3071), .D(n3145), .Q(
        \bank_register[24][1] ) );
  DLH_X1 \bank_register_reg[24][0]  ( .G(n3070), .D(n3142), .Q(
        \bank_register[24][0] ) );
  DLH_X1 \bank_register_reg[25][31]  ( .G(n3069), .D(n3235), .Q(
        \bank_register[25][31] ) );
  DLH_X1 \bank_register_reg[25][30]  ( .G(n3069), .D(n3232), .Q(
        \bank_register[25][30] ) );
  DLH_X1 \bank_register_reg[25][29]  ( .G(n3067), .D(n3229), .Q(
        \bank_register[25][29] ) );
  DLH_X1 \bank_register_reg[25][28]  ( .G(n3067), .D(n3226), .Q(
        \bank_register[25][28] ) );
  DLH_X1 \bank_register_reg[25][27]  ( .G(n3067), .D(n3223), .Q(
        \bank_register[25][27] ) );
  DLH_X1 \bank_register_reg[25][26]  ( .G(n3067), .D(n3220), .Q(
        \bank_register[25][26] ) );
  DLH_X1 \bank_register_reg[25][25]  ( .G(n3067), .D(n3217), .Q(
        \bank_register[25][25] ) );
  DLH_X1 \bank_register_reg[25][24]  ( .G(n3067), .D(n3214), .Q(
        \bank_register[25][24] ) );
  DLH_X1 \bank_register_reg[25][23]  ( .G(n3067), .D(n3211), .Q(
        \bank_register[25][23] ) );
  DLH_X1 \bank_register_reg[25][22]  ( .G(n3067), .D(n3208), .Q(
        \bank_register[25][22] ) );
  DLH_X1 \bank_register_reg[25][21]  ( .G(n3067), .D(n3205), .Q(
        \bank_register[25][21] ) );
  DLH_X1 \bank_register_reg[25][20]  ( .G(n3067), .D(n3202), .Q(
        \bank_register[25][20] ) );
  DLH_X1 \bank_register_reg[25][19]  ( .G(n3068), .D(n3199), .Q(
        \bank_register[25][19] ) );
  DLH_X1 \bank_register_reg[25][18]  ( .G(n3068), .D(n3196), .Q(
        \bank_register[25][18] ) );
  DLH_X1 \bank_register_reg[25][17]  ( .G(n3069), .D(n3193), .Q(
        \bank_register[25][17] ) );
  DLH_X1 \bank_register_reg[25][16]  ( .G(n3069), .D(n3190), .Q(
        \bank_register[25][16] ) );
  DLH_X1 \bank_register_reg[25][15]  ( .G(n3069), .D(n3187), .Q(
        \bank_register[25][15] ) );
  DLH_X1 \bank_register_reg[25][14]  ( .G(n3069), .D(n3184), .Q(
        \bank_register[25][14] ) );
  DLH_X1 \bank_register_reg[25][13]  ( .G(n3069), .D(n3181), .Q(
        \bank_register[25][13] ) );
  DLH_X1 \bank_register_reg[25][12]  ( .G(n3069), .D(n3178), .Q(
        \bank_register[25][12] ) );
  DLH_X1 \bank_register_reg[25][11]  ( .G(n3069), .D(n3175), .Q(
        \bank_register[25][11] ) );
  DLH_X1 \bank_register_reg[25][10]  ( .G(n3069), .D(n3172), .Q(
        \bank_register[25][10] ) );
  DLH_X1 \bank_register_reg[25][9]  ( .G(n3068), .D(n3169), .Q(
        \bank_register[25][9] ) );
  DLH_X1 \bank_register_reg[25][8]  ( .G(n3068), .D(n3166), .Q(
        \bank_register[25][8] ) );
  DLH_X1 \bank_register_reg[25][7]  ( .G(n3068), .D(n3163), .Q(
        \bank_register[25][7] ) );
  DLH_X1 \bank_register_reg[25][6]  ( .G(n3068), .D(n3160), .Q(
        \bank_register[25][6] ) );
  DLH_X1 \bank_register_reg[25][5]  ( .G(n3068), .D(n3157), .Q(
        \bank_register[25][5] ) );
  DLH_X1 \bank_register_reg[25][4]  ( .G(n3068), .D(n3154), .Q(
        \bank_register[25][4] ) );
  DLH_X1 \bank_register_reg[25][3]  ( .G(n3068), .D(n3151), .Q(
        \bank_register[25][3] ) );
  DLH_X1 \bank_register_reg[25][2]  ( .G(n3068), .D(n3148), .Q(
        \bank_register[25][2] ) );
  DLH_X1 \bank_register_reg[25][1]  ( .G(n3068), .D(n3145), .Q(
        \bank_register[25][1] ) );
  DLH_X1 \bank_register_reg[25][0]  ( .G(n3067), .D(n3142), .Q(
        \bank_register[25][0] ) );
  DLH_X1 \bank_register_reg[26][31]  ( .G(n3066), .D(n3235), .Q(
        \bank_register[26][31] ) );
  DLH_X1 \bank_register_reg[26][30]  ( .G(n3066), .D(n3232), .Q(
        \bank_register[26][30] ) );
  DLH_X1 \bank_register_reg[26][29]  ( .G(n3064), .D(n3229), .Q(
        \bank_register[26][29] ) );
  DLH_X1 \bank_register_reg[26][28]  ( .G(n3064), .D(n3226), .Q(
        \bank_register[26][28] ) );
  DLH_X1 \bank_register_reg[26][27]  ( .G(n3064), .D(n3223), .Q(
        \bank_register[26][27] ) );
  DLH_X1 \bank_register_reg[26][26]  ( .G(n3064), .D(n3220), .Q(
        \bank_register[26][26] ) );
  DLH_X1 \bank_register_reg[26][25]  ( .G(n3064), .D(n3217), .Q(
        \bank_register[26][25] ) );
  DLH_X1 \bank_register_reg[26][24]  ( .G(n3064), .D(n3214), .Q(
        \bank_register[26][24] ) );
  DLH_X1 \bank_register_reg[26][23]  ( .G(n3064), .D(n3211), .Q(
        \bank_register[26][23] ) );
  DLH_X1 \bank_register_reg[26][22]  ( .G(n3064), .D(n3208), .Q(
        \bank_register[26][22] ) );
  DLH_X1 \bank_register_reg[26][21]  ( .G(n3064), .D(n3205), .Q(
        \bank_register[26][21] ) );
  DLH_X1 \bank_register_reg[26][20]  ( .G(n3064), .D(n3202), .Q(
        \bank_register[26][20] ) );
  DLH_X1 \bank_register_reg[26][19]  ( .G(n3065), .D(n3199), .Q(
        \bank_register[26][19] ) );
  DLH_X1 \bank_register_reg[26][18]  ( .G(n3065), .D(n3196), .Q(
        \bank_register[26][18] ) );
  DLH_X1 \bank_register_reg[26][17]  ( .G(n3066), .D(n3193), .Q(
        \bank_register[26][17] ) );
  DLH_X1 \bank_register_reg[26][16]  ( .G(n3066), .D(n3190), .Q(
        \bank_register[26][16] ) );
  DLH_X1 \bank_register_reg[26][15]  ( .G(n3066), .D(n3187), .Q(
        \bank_register[26][15] ) );
  DLH_X1 \bank_register_reg[26][14]  ( .G(n3066), .D(n3184), .Q(
        \bank_register[26][14] ) );
  DLH_X1 \bank_register_reg[26][13]  ( .G(n3066), .D(n3181), .Q(
        \bank_register[26][13] ) );
  DLH_X1 \bank_register_reg[26][12]  ( .G(n3066), .D(n3178), .Q(
        \bank_register[26][12] ) );
  DLH_X1 \bank_register_reg[26][11]  ( .G(n3066), .D(n3175), .Q(
        \bank_register[26][11] ) );
  DLH_X1 \bank_register_reg[26][10]  ( .G(n3066), .D(n3172), .Q(
        \bank_register[26][10] ) );
  DLH_X1 \bank_register_reg[26][9]  ( .G(n3065), .D(n3169), .Q(
        \bank_register[26][9] ) );
  DLH_X1 \bank_register_reg[26][8]  ( .G(n3065), .D(n3166), .Q(
        \bank_register[26][8] ) );
  DLH_X1 \bank_register_reg[26][7]  ( .G(n3065), .D(n3163), .Q(
        \bank_register[26][7] ) );
  DLH_X1 \bank_register_reg[26][6]  ( .G(n3065), .D(n3160), .Q(
        \bank_register[26][6] ) );
  DLH_X1 \bank_register_reg[26][5]  ( .G(n3065), .D(n3157), .Q(
        \bank_register[26][5] ) );
  DLH_X1 \bank_register_reg[26][4]  ( .G(n3065), .D(n3154), .Q(
        \bank_register[26][4] ) );
  DLH_X1 \bank_register_reg[26][3]  ( .G(n3065), .D(n3151), .Q(
        \bank_register[26][3] ) );
  DLH_X1 \bank_register_reg[26][2]  ( .G(n3065), .D(n3148), .Q(
        \bank_register[26][2] ) );
  DLH_X1 \bank_register_reg[26][1]  ( .G(n3065), .D(n3145), .Q(
        \bank_register[26][1] ) );
  DLH_X1 \bank_register_reg[26][0]  ( .G(n3064), .D(n3142), .Q(
        \bank_register[26][0] ) );
  DLH_X1 \bank_register_reg[27][31]  ( .G(n3063), .D(n3235), .Q(
        \bank_register[27][31] ) );
  DLH_X1 \bank_register_reg[27][30]  ( .G(n3063), .D(n3232), .Q(
        \bank_register[27][30] ) );
  DLH_X1 \bank_register_reg[27][29]  ( .G(n3061), .D(n3229), .Q(
        \bank_register[27][29] ) );
  DLH_X1 \bank_register_reg[27][28]  ( .G(n3061), .D(n3226), .Q(
        \bank_register[27][28] ) );
  DLH_X1 \bank_register_reg[27][27]  ( .G(n3061), .D(n3223), .Q(
        \bank_register[27][27] ) );
  DLH_X1 \bank_register_reg[27][26]  ( .G(n3061), .D(n3220), .Q(
        \bank_register[27][26] ) );
  DLH_X1 \bank_register_reg[27][25]  ( .G(n3061), .D(n3217), .Q(
        \bank_register[27][25] ) );
  DLH_X1 \bank_register_reg[27][24]  ( .G(n3061), .D(n3214), .Q(
        \bank_register[27][24] ) );
  DLH_X1 \bank_register_reg[27][23]  ( .G(n3061), .D(n3211), .Q(
        \bank_register[27][23] ) );
  DLH_X1 \bank_register_reg[27][22]  ( .G(n3061), .D(n3208), .Q(
        \bank_register[27][22] ) );
  DLH_X1 \bank_register_reg[27][21]  ( .G(n3061), .D(n3205), .Q(
        \bank_register[27][21] ) );
  DLH_X1 \bank_register_reg[27][20]  ( .G(n3061), .D(n3202), .Q(
        \bank_register[27][20] ) );
  DLH_X1 \bank_register_reg[27][19]  ( .G(n3062), .D(n3199), .Q(
        \bank_register[27][19] ) );
  DLH_X1 \bank_register_reg[27][18]  ( .G(n3062), .D(n3196), .Q(
        \bank_register[27][18] ) );
  DLH_X1 \bank_register_reg[27][17]  ( .G(n3063), .D(n3193), .Q(
        \bank_register[27][17] ) );
  DLH_X1 \bank_register_reg[27][16]  ( .G(n3063), .D(n3190), .Q(
        \bank_register[27][16] ) );
  DLH_X1 \bank_register_reg[27][15]  ( .G(n3063), .D(n3187), .Q(
        \bank_register[27][15] ) );
  DLH_X1 \bank_register_reg[27][14]  ( .G(n3063), .D(n3184), .Q(
        \bank_register[27][14] ) );
  DLH_X1 \bank_register_reg[27][13]  ( .G(n3063), .D(n3181), .Q(
        \bank_register[27][13] ) );
  DLH_X1 \bank_register_reg[27][12]  ( .G(n3063), .D(n3178), .Q(
        \bank_register[27][12] ) );
  DLH_X1 \bank_register_reg[27][11]  ( .G(n3063), .D(n3175), .Q(
        \bank_register[27][11] ) );
  DLH_X1 \bank_register_reg[27][10]  ( .G(n3063), .D(n3172), .Q(
        \bank_register[27][10] ) );
  DLH_X1 \bank_register_reg[27][9]  ( .G(n3062), .D(n3169), .Q(
        \bank_register[27][9] ) );
  DLH_X1 \bank_register_reg[27][8]  ( .G(n3062), .D(n3166), .Q(
        \bank_register[27][8] ) );
  DLH_X1 \bank_register_reg[27][7]  ( .G(n3062), .D(n3163), .Q(
        \bank_register[27][7] ) );
  DLH_X1 \bank_register_reg[27][6]  ( .G(n3062), .D(n3160), .Q(
        \bank_register[27][6] ) );
  DLH_X1 \bank_register_reg[27][5]  ( .G(n3062), .D(n3157), .Q(
        \bank_register[27][5] ) );
  DLH_X1 \bank_register_reg[27][4]  ( .G(n3062), .D(n3154), .Q(
        \bank_register[27][4] ) );
  DLH_X1 \bank_register_reg[27][3]  ( .G(n3062), .D(n3151), .Q(
        \bank_register[27][3] ) );
  DLH_X1 \bank_register_reg[27][2]  ( .G(n3062), .D(n3148), .Q(
        \bank_register[27][2] ) );
  DLH_X1 \bank_register_reg[27][1]  ( .G(n3062), .D(n3145), .Q(
        \bank_register[27][1] ) );
  DLH_X1 \bank_register_reg[27][0]  ( .G(n3061), .D(n3142), .Q(
        \bank_register[27][0] ) );
  DLH_X1 \bank_register_reg[28][31]  ( .G(n3060), .D(n3235), .Q(
        \bank_register[28][31] ) );
  DLH_X1 \bank_register_reg[28][30]  ( .G(n3060), .D(n3232), .Q(
        \bank_register[28][30] ) );
  DLH_X1 \bank_register_reg[28][29]  ( .G(n3058), .D(n3229), .Q(
        \bank_register[28][29] ) );
  DLH_X1 \bank_register_reg[28][28]  ( .G(n3058), .D(n3226), .Q(
        \bank_register[28][28] ) );
  DLH_X1 \bank_register_reg[28][27]  ( .G(n3058), .D(n3223), .Q(
        \bank_register[28][27] ) );
  DLH_X1 \bank_register_reg[28][26]  ( .G(n3058), .D(n3220), .Q(
        \bank_register[28][26] ) );
  DLH_X1 \bank_register_reg[28][25]  ( .G(n3058), .D(n3217), .Q(
        \bank_register[28][25] ) );
  DLH_X1 \bank_register_reg[28][24]  ( .G(n3058), .D(n3214), .Q(
        \bank_register[28][24] ) );
  DLH_X1 \bank_register_reg[28][23]  ( .G(n3058), .D(n3211), .Q(
        \bank_register[28][23] ) );
  DLH_X1 \bank_register_reg[28][22]  ( .G(n3058), .D(n3208), .Q(
        \bank_register[28][22] ) );
  DLH_X1 \bank_register_reg[28][21]  ( .G(n3058), .D(n3205), .Q(
        \bank_register[28][21] ) );
  DLH_X1 \bank_register_reg[28][20]  ( .G(n3058), .D(n3202), .Q(
        \bank_register[28][20] ) );
  DLH_X1 \bank_register_reg[28][19]  ( .G(n3059), .D(n3199), .Q(
        \bank_register[28][19] ) );
  DLH_X1 \bank_register_reg[28][18]  ( .G(n3059), .D(n3196), .Q(
        \bank_register[28][18] ) );
  DLH_X1 \bank_register_reg[28][17]  ( .G(n3060), .D(n3193), .Q(
        \bank_register[28][17] ) );
  DLH_X1 \bank_register_reg[28][16]  ( .G(n3060), .D(n3190), .Q(
        \bank_register[28][16] ) );
  DLH_X1 \bank_register_reg[28][15]  ( .G(n3060), .D(n3187), .Q(
        \bank_register[28][15] ) );
  DLH_X1 \bank_register_reg[28][14]  ( .G(n3060), .D(n3184), .Q(
        \bank_register[28][14] ) );
  DLH_X1 \bank_register_reg[28][13]  ( .G(n3060), .D(n3181), .Q(
        \bank_register[28][13] ) );
  DLH_X1 \bank_register_reg[28][12]  ( .G(n3060), .D(n3178), .Q(
        \bank_register[28][12] ) );
  DLH_X1 \bank_register_reg[28][11]  ( .G(n3060), .D(n3175), .Q(
        \bank_register[28][11] ) );
  DLH_X1 \bank_register_reg[28][10]  ( .G(n3060), .D(n3172), .Q(
        \bank_register[28][10] ) );
  DLH_X1 \bank_register_reg[28][9]  ( .G(n3059), .D(n3169), .Q(
        \bank_register[28][9] ) );
  DLH_X1 \bank_register_reg[28][8]  ( .G(n3059), .D(n3166), .Q(
        \bank_register[28][8] ) );
  DLH_X1 \bank_register_reg[28][7]  ( .G(n3059), .D(n3163), .Q(
        \bank_register[28][7] ) );
  DLH_X1 \bank_register_reg[28][6]  ( .G(n3059), .D(n3160), .Q(
        \bank_register[28][6] ) );
  DLH_X1 \bank_register_reg[28][5]  ( .G(n3059), .D(n3157), .Q(
        \bank_register[28][5] ) );
  DLH_X1 \bank_register_reg[28][4]  ( .G(n3059), .D(n3154), .Q(
        \bank_register[28][4] ) );
  DLH_X1 \bank_register_reg[28][3]  ( .G(n3059), .D(n3151), .Q(
        \bank_register[28][3] ) );
  DLH_X1 \bank_register_reg[28][2]  ( .G(n3059), .D(n3148), .Q(
        \bank_register[28][2] ) );
  DLH_X1 \bank_register_reg[28][1]  ( .G(n3059), .D(n3145), .Q(
        \bank_register[28][1] ) );
  DLH_X1 \bank_register_reg[28][0]  ( .G(n3058), .D(n3142), .Q(
        \bank_register[28][0] ) );
  DLH_X1 \bank_register_reg[29][31]  ( .G(n3057), .D(n3235), .Q(
        \bank_register[29][31] ) );
  DLH_X1 \bank_register_reg[29][30]  ( .G(n3057), .D(n3232), .Q(
        \bank_register[29][30] ) );
  DLH_X1 \bank_register_reg[29][29]  ( .G(n3055), .D(n3229), .Q(
        \bank_register[29][29] ) );
  DLH_X1 \bank_register_reg[29][28]  ( .G(n3055), .D(n3226), .Q(
        \bank_register[29][28] ) );
  DLH_X1 \bank_register_reg[29][27]  ( .G(n3055), .D(n3223), .Q(
        \bank_register[29][27] ) );
  DLH_X1 \bank_register_reg[29][26]  ( .G(n3055), .D(n3220), .Q(
        \bank_register[29][26] ) );
  DLH_X1 \bank_register_reg[29][25]  ( .G(n3055), .D(n3217), .Q(
        \bank_register[29][25] ) );
  DLH_X1 \bank_register_reg[29][24]  ( .G(n3055), .D(n3214), .Q(
        \bank_register[29][24] ) );
  DLH_X1 \bank_register_reg[29][23]  ( .G(n3055), .D(n3211), .Q(
        \bank_register[29][23] ) );
  DLH_X1 \bank_register_reg[29][22]  ( .G(n3055), .D(n3208), .Q(
        \bank_register[29][22] ) );
  DLH_X1 \bank_register_reg[29][21]  ( .G(n3055), .D(n3205), .Q(
        \bank_register[29][21] ) );
  DLH_X1 \bank_register_reg[29][20]  ( .G(n3055), .D(n3202), .Q(
        \bank_register[29][20] ) );
  DLH_X1 \bank_register_reg[29][19]  ( .G(n3056), .D(n3199), .Q(
        \bank_register[29][19] ) );
  DLH_X1 \bank_register_reg[29][18]  ( .G(n3056), .D(n3196), .Q(
        \bank_register[29][18] ) );
  DLH_X1 \bank_register_reg[29][17]  ( .G(n3057), .D(n3193), .Q(
        \bank_register[29][17] ) );
  DLH_X1 \bank_register_reg[29][16]  ( .G(n3057), .D(n3190), .Q(
        \bank_register[29][16] ) );
  DLH_X1 \bank_register_reg[29][15]  ( .G(n3057), .D(n3187), .Q(
        \bank_register[29][15] ) );
  DLH_X1 \bank_register_reg[29][14]  ( .G(n3057), .D(n3184), .Q(
        \bank_register[29][14] ) );
  DLH_X1 \bank_register_reg[29][13]  ( .G(n3057), .D(n3181), .Q(
        \bank_register[29][13] ) );
  DLH_X1 \bank_register_reg[29][12]  ( .G(n3057), .D(n3178), .Q(
        \bank_register[29][12] ) );
  DLH_X1 \bank_register_reg[29][11]  ( .G(n3057), .D(n3175), .Q(
        \bank_register[29][11] ) );
  DLH_X1 \bank_register_reg[29][10]  ( .G(n3057), .D(n3172), .Q(
        \bank_register[29][10] ) );
  DLH_X1 \bank_register_reg[29][9]  ( .G(n3056), .D(n3169), .Q(
        \bank_register[29][9] ) );
  DLH_X1 \bank_register_reg[29][8]  ( .G(n3056), .D(n3166), .Q(
        \bank_register[29][8] ) );
  DLH_X1 \bank_register_reg[29][7]  ( .G(n3056), .D(n3163), .Q(
        \bank_register[29][7] ) );
  DLH_X1 \bank_register_reg[29][6]  ( .G(n3056), .D(n3160), .Q(
        \bank_register[29][6] ) );
  DLH_X1 \bank_register_reg[29][5]  ( .G(n3056), .D(n3157), .Q(
        \bank_register[29][5] ) );
  DLH_X1 \bank_register_reg[29][4]  ( .G(n3056), .D(n3154), .Q(
        \bank_register[29][4] ) );
  DLH_X1 \bank_register_reg[29][3]  ( .G(n3056), .D(n3151), .Q(
        \bank_register[29][3] ) );
  DLH_X1 \bank_register_reg[29][2]  ( .G(n3056), .D(n3148), .Q(
        \bank_register[29][2] ) );
  DLH_X1 \bank_register_reg[29][1]  ( .G(n3056), .D(n3145), .Q(
        \bank_register[29][1] ) );
  DLH_X1 \bank_register_reg[29][0]  ( .G(n3055), .D(n3142), .Q(
        \bank_register[29][0] ) );
  DLH_X1 \bank_register_reg[30][31]  ( .G(n3054), .D(n3235), .Q(
        \bank_register[30][31] ) );
  DLH_X1 \bank_register_reg[30][30]  ( .G(n3054), .D(n3232), .Q(
        \bank_register[30][30] ) );
  DLH_X1 \bank_register_reg[30][29]  ( .G(n3052), .D(n3229), .Q(
        \bank_register[30][29] ) );
  DLH_X1 \bank_register_reg[30][28]  ( .G(n3052), .D(n3226), .Q(
        \bank_register[30][28] ) );
  DLH_X1 \bank_register_reg[30][27]  ( .G(n3052), .D(n3223), .Q(
        \bank_register[30][27] ) );
  DLH_X1 \bank_register_reg[30][26]  ( .G(n3052), .D(n3220), .Q(
        \bank_register[30][26] ) );
  DLH_X1 \bank_register_reg[30][25]  ( .G(n3052), .D(n3217), .Q(
        \bank_register[30][25] ) );
  DLH_X1 \bank_register_reg[30][24]  ( .G(n3052), .D(n3214), .Q(
        \bank_register[30][24] ) );
  DLH_X1 \bank_register_reg[30][23]  ( .G(n3052), .D(n3211), .Q(
        \bank_register[30][23] ) );
  DLH_X1 \bank_register_reg[30][22]  ( .G(n3052), .D(n3208), .Q(
        \bank_register[30][22] ) );
  DLH_X1 \bank_register_reg[30][21]  ( .G(n3052), .D(n3205), .Q(
        \bank_register[30][21] ) );
  DLH_X1 \bank_register_reg[30][20]  ( .G(n3052), .D(n3202), .Q(
        \bank_register[30][20] ) );
  DLH_X1 \bank_register_reg[30][19]  ( .G(n3053), .D(n3199), .Q(
        \bank_register[30][19] ) );
  DLH_X1 \bank_register_reg[30][18]  ( .G(n3053), .D(n3196), .Q(
        \bank_register[30][18] ) );
  DLH_X1 \bank_register_reg[30][17]  ( .G(n3054), .D(n3193), .Q(
        \bank_register[30][17] ) );
  DLH_X1 \bank_register_reg[30][16]  ( .G(n3054), .D(n3190), .Q(
        \bank_register[30][16] ) );
  DLH_X1 \bank_register_reg[30][15]  ( .G(n3054), .D(n3187), .Q(
        \bank_register[30][15] ) );
  DLH_X1 \bank_register_reg[30][14]  ( .G(n3054), .D(n3184), .Q(
        \bank_register[30][14] ) );
  DLH_X1 \bank_register_reg[30][13]  ( .G(n3054), .D(n3181), .Q(
        \bank_register[30][13] ) );
  DLH_X1 \bank_register_reg[30][12]  ( .G(n3054), .D(n3178), .Q(
        \bank_register[30][12] ) );
  DLH_X1 \bank_register_reg[30][11]  ( .G(n3054), .D(n3175), .Q(
        \bank_register[30][11] ) );
  DLH_X1 \bank_register_reg[30][10]  ( .G(n3054), .D(n3172), .Q(
        \bank_register[30][10] ) );
  DLH_X1 \bank_register_reg[30][9]  ( .G(n3053), .D(n3169), .Q(
        \bank_register[30][9] ) );
  DLH_X1 \bank_register_reg[30][8]  ( .G(n3053), .D(n3166), .Q(
        \bank_register[30][8] ) );
  DLH_X1 \bank_register_reg[30][7]  ( .G(n3053), .D(n3163), .Q(
        \bank_register[30][7] ) );
  DLH_X1 \bank_register_reg[30][6]  ( .G(n3053), .D(n3160), .Q(
        \bank_register[30][6] ) );
  DLH_X1 \bank_register_reg[30][5]  ( .G(n3053), .D(n3157), .Q(
        \bank_register[30][5] ) );
  DLH_X1 \bank_register_reg[30][4]  ( .G(n3053), .D(n3154), .Q(
        \bank_register[30][4] ) );
  DLH_X1 \bank_register_reg[30][3]  ( .G(n3053), .D(n3151), .Q(
        \bank_register[30][3] ) );
  DLH_X1 \bank_register_reg[30][2]  ( .G(n3053), .D(n3148), .Q(
        \bank_register[30][2] ) );
  DLH_X1 \bank_register_reg[30][1]  ( .G(n3053), .D(n3145), .Q(
        \bank_register[30][1] ) );
  DLH_X1 \bank_register_reg[30][0]  ( .G(n3052), .D(n3142), .Q(
        \bank_register[30][0] ) );
  DLH_X1 \bank_register_reg[31][31]  ( .G(n3051), .D(n3236), .Q(
        \bank_register[31][31] ) );
  DLH_X1 \bank_register_reg[31][30]  ( .G(n3051), .D(n3233), .Q(
        \bank_register[31][30] ) );
  DLH_X1 \bank_register_reg[31][29]  ( .G(n3049), .D(n3230), .Q(
        \bank_register[31][29] ) );
  DLH_X1 \bank_register_reg[31][28]  ( .G(n3049), .D(n3227), .Q(
        \bank_register[31][28] ) );
  DLH_X1 \bank_register_reg[31][27]  ( .G(n3049), .D(n3224), .Q(
        \bank_register[31][27] ) );
  DLH_X1 \bank_register_reg[31][26]  ( .G(n3049), .D(n3221), .Q(
        \bank_register[31][26] ) );
  DLH_X1 \bank_register_reg[31][25]  ( .G(n3049), .D(n3218), .Q(
        \bank_register[31][25] ) );
  DLH_X1 \bank_register_reg[31][24]  ( .G(n3049), .D(n3215), .Q(
        \bank_register[31][24] ) );
  DLH_X1 \bank_register_reg[31][23]  ( .G(n3049), .D(n3212), .Q(
        \bank_register[31][23] ) );
  DLH_X1 \bank_register_reg[31][22]  ( .G(n3049), .D(n3209), .Q(
        \bank_register[31][22] ) );
  DLH_X1 \bank_register_reg[31][21]  ( .G(n3049), .D(n3206), .Q(
        \bank_register[31][21] ) );
  DLH_X1 \bank_register_reg[31][20]  ( .G(n3049), .D(n3203), .Q(
        \bank_register[31][20] ) );
  DLH_X1 \bank_register_reg[31][19]  ( .G(n3050), .D(n3200), .Q(
        \bank_register[31][19] ) );
  DLH_X1 \bank_register_reg[31][18]  ( .G(n3050), .D(n3197), .Q(
        \bank_register[31][18] ) );
  DLH_X1 \bank_register_reg[31][17]  ( .G(n3051), .D(n3194), .Q(
        \bank_register[31][17] ) );
  DLH_X1 \bank_register_reg[31][16]  ( .G(n3051), .D(n3191), .Q(
        \bank_register[31][16] ) );
  DLH_X1 \bank_register_reg[31][15]  ( .G(n3051), .D(n3188), .Q(
        \bank_register[31][15] ) );
  DLH_X1 \bank_register_reg[31][14]  ( .G(n3051), .D(n3185), .Q(
        \bank_register[31][14] ) );
  DLH_X1 \bank_register_reg[31][13]  ( .G(n3051), .D(n3182), .Q(
        \bank_register[31][13] ) );
  DLH_X1 \bank_register_reg[31][12]  ( .G(n3051), .D(n3179), .Q(
        \bank_register[31][12] ) );
  DLH_X1 \bank_register_reg[31][11]  ( .G(n3051), .D(n3176), .Q(
        \bank_register[31][11] ) );
  DLH_X1 \bank_register_reg[31][10]  ( .G(n3051), .D(n3173), .Q(
        \bank_register[31][10] ) );
  DLH_X1 \bank_register_reg[31][9]  ( .G(n3050), .D(n3170), .Q(
        \bank_register[31][9] ) );
  DLH_X1 \bank_register_reg[31][8]  ( .G(n3050), .D(n3167), .Q(
        \bank_register[31][8] ) );
  DLH_X1 \bank_register_reg[31][7]  ( .G(n3050), .D(n3164), .Q(
        \bank_register[31][7] ) );
  DLH_X1 \bank_register_reg[31][6]  ( .G(n3050), .D(n3161), .Q(
        \bank_register[31][6] ) );
  DLH_X1 \bank_register_reg[31][5]  ( .G(n3050), .D(n3158), .Q(
        \bank_register[31][5] ) );
  DLH_X1 \bank_register_reg[31][4]  ( .G(n3050), .D(n3155), .Q(
        \bank_register[31][4] ) );
  DLH_X1 \bank_register_reg[31][3]  ( .G(n3050), .D(n3152), .Q(
        \bank_register[31][3] ) );
  DLH_X1 \bank_register_reg[31][2]  ( .G(n3050), .D(n3149), .Q(
        \bank_register[31][2] ) );
  DLH_X1 \bank_register_reg[31][1]  ( .G(n3050), .D(n3146), .Q(
        \bank_register[31][1] ) );
  DLH_X1 \bank_register_reg[31][0]  ( .G(n3049), .D(n3143), .Q(
        \bank_register[31][0] ) );
  NAND3_X1 U2179 ( .A1(write_address[3]), .A2(reg_write), .A3(write_address[4]), .ZN(n662) );
  NAND3_X1 U2180 ( .A1(reg_write), .A2(n673), .A3(write_address[4]), .ZN(n672)
         );
  NAND3_X1 U2181 ( .A1(reg_write), .A2(n675), .A3(write_address[3]), .ZN(n674)
         );
  NAND3_X1 U2182 ( .A1(n676), .A2(n677), .A3(n678), .ZN(n671) );
  NAND3_X1 U2183 ( .A1(write_address[1]), .A2(write_address[0]), .A3(
        write_address[2]), .ZN(n663) );
  NAND3_X1 U2184 ( .A1(write_address[1]), .A2(n678), .A3(write_address[2]), 
        .ZN(n665) );
  NAND3_X1 U2185 ( .A1(write_address[0]), .A2(n676), .A3(write_address[2]), 
        .ZN(n666) );
  NAND3_X1 U2186 ( .A1(n678), .A2(n676), .A3(write_address[2]), .ZN(n667) );
  NAND3_X1 U2187 ( .A1(write_address[0]), .A2(n677), .A3(write_address[1]), 
        .ZN(n668) );
  NAND3_X1 U2188 ( .A1(n678), .A2(n677), .A3(write_address[1]), .ZN(n669) );
  NAND3_X1 U2189 ( .A1(n673), .A2(n675), .A3(reg_write), .ZN(n679) );
  NAND3_X1 U2190 ( .A1(n676), .A2(n677), .A3(write_address[0]), .ZN(n670) );
  XOR2_X1 U2191 ( .A(write_address[4]), .B(read_address_2[4]), .Z(n1887) );
  XOR2_X1 U2192 ( .A(write_address[2]), .B(read_address_2[2]), .Z(n1886) );
  XOR2_X1 U2193 ( .A(n678), .B(read_address_2[0]), .Z(n1882) );
  XOR2_X1 U2194 ( .A(n1879), .B(write_address[1]), .Z(n1881) );
  XOR2_X1 U2195 ( .A(n1888), .B(write_address[3]), .Z(n1880) );
  NAND3_X1 U2196 ( .A1(n1888), .A2(n1895), .A3(n1896), .ZN(n714) );
  NAND3_X1 U2197 ( .A1(n1888), .A2(n1895), .A3(read_address_2[2]), .ZN(n712)
         );
  NAND3_X1 U2198 ( .A1(n2785), .A2(n2786), .A3(n2787), .ZN(n1911) );
  NAND3_X1 U2199 ( .A1(n2785), .A2(n2786), .A3(read_address_1[2]), .ZN(n1912)
         );
  XOR2_X1 U2200 ( .A(write_address[4]), .B(read_address_1[4]), .Z(n2799) );
  XOR2_X1 U2201 ( .A(write_address[2]), .B(read_address_1[2]), .Z(n2798) );
  XOR2_X1 U2202 ( .A(n678), .B(n3240), .Z(n2796) );
  XOR2_X1 U2203 ( .A(read_address_1[1]), .B(n676), .Z(n2795) );
  XOR2_X1 U2204 ( .A(n2785), .B(write_address[3]), .Z(n2794) );
  BUF_X1 U3 ( .A(n2997), .Z(n3001) );
  BUF_X1 U4 ( .A(n2997), .Z(n3000) );
  BUF_X1 U5 ( .A(n2997), .Z(n3002) );
  BUF_X1 U6 ( .A(n2998), .Z(n3003) );
  BUF_X1 U7 ( .A(n2998), .Z(n3004) );
  BUF_X1 U8 ( .A(n2998), .Z(n3005) );
  BUF_X1 U9 ( .A(n2999), .Z(n3007) );
  BUF_X1 U10 ( .A(n2999), .Z(n3006) );
  BUF_X1 U11 ( .A(n683), .Z(n3036) );
  BUF_X1 U12 ( .A(n683), .Z(n3037) );
  BUF_X1 U13 ( .A(n683), .Z(n3038) );
  BUF_X1 U14 ( .A(n1934), .Z(n2811) );
  BUF_X1 U15 ( .A(n1945), .Z(n2802) );
  BUF_X1 U16 ( .A(n1934), .Z(n2812) );
  BUF_X1 U17 ( .A(n1945), .Z(n2803) );
  BUF_X1 U18 ( .A(n1946), .Z(n2767) );
  BUF_X1 U19 ( .A(n1946), .Z(n2800) );
  BUF_X1 U20 ( .A(n2986), .Z(n2990) );
  BUF_X1 U21 ( .A(n2942), .Z(n2946) );
  BUF_X1 U22 ( .A(n2986), .Z(n2989) );
  BUF_X1 U23 ( .A(n2942), .Z(n2945) );
  BUF_X1 U24 ( .A(n2987), .Z(n2992) );
  BUF_X1 U25 ( .A(n2943), .Z(n2948) );
  BUF_X1 U26 ( .A(n2987), .Z(n2993) );
  BUF_X1 U27 ( .A(n2943), .Z(n2949) );
  BUF_X1 U28 ( .A(n2943), .Z(n2950) );
  BUF_X1 U29 ( .A(n2987), .Z(n2994) );
  BUF_X1 U30 ( .A(n692), .Z(n3027) );
  BUF_X1 U31 ( .A(n694), .Z(n3021) );
  BUF_X1 U32 ( .A(n692), .Z(n3028) );
  BUF_X1 U33 ( .A(n694), .Z(n3022) );
  BUF_X1 U34 ( .A(n2988), .Z(n2995) );
  BUF_X1 U35 ( .A(n2944), .Z(n2951) );
  BUF_X1 U36 ( .A(n3008), .Z(n3009) );
  BUF_X1 U37 ( .A(n3008), .Z(n3010) );
  BUF_X1 U38 ( .A(n2904), .Z(n2911) );
  BUF_X1 U39 ( .A(n2860), .Z(n2867) );
  BUF_X1 U40 ( .A(n2904), .Z(n2910) );
  BUF_X1 U41 ( .A(n2860), .Z(n2866) );
  BUF_X1 U42 ( .A(n2904), .Z(n2909) );
  BUF_X1 U43 ( .A(n2860), .Z(n2865) );
  BUF_X1 U44 ( .A(n2861), .Z(n2868) );
  BUF_X1 U45 ( .A(n2905), .Z(n2912) );
  BUF_X1 U46 ( .A(n693), .Z(n3024) );
  BUF_X1 U47 ( .A(n693), .Z(n3025) );
  BUF_X1 U48 ( .A(n2848), .Z(n2851) );
  BUF_X1 U49 ( .A(n2848), .Z(n2852) );
  BUF_X1 U50 ( .A(n2986), .Z(n2991) );
  BUF_X1 U51 ( .A(n2942), .Z(n2947) );
  BUF_X1 U52 ( .A(n2848), .Z(n2853) );
  BUF_X1 U53 ( .A(n2859), .Z(n2862) );
  BUF_X1 U54 ( .A(n2903), .Z(n2906) );
  BUF_X1 U55 ( .A(n2859), .Z(n2863) );
  BUF_X1 U56 ( .A(n2903), .Z(n2907) );
  BUF_X1 U57 ( .A(n2859), .Z(n2864) );
  BUF_X1 U58 ( .A(n2903), .Z(n2908) );
  BUF_X1 U59 ( .A(n2849), .Z(n2856) );
  BUF_X1 U60 ( .A(n2849), .Z(n2855) );
  BUF_X1 U61 ( .A(n2849), .Z(n2854) );
  BUF_X1 U62 ( .A(n2850), .Z(n2858) );
  BUF_X1 U63 ( .A(n2850), .Z(n2857) );
  BUF_X1 U64 ( .A(n2837), .Z(n2840) );
  BUF_X1 U65 ( .A(n2837), .Z(n2841) );
  BUF_X1 U66 ( .A(n2837), .Z(n2842) );
  BUF_X1 U67 ( .A(n2964), .Z(n2967) );
  BUF_X1 U68 ( .A(n2920), .Z(n2923) );
  BUF_X1 U69 ( .A(n2920), .Z(n2924) );
  BUF_X1 U70 ( .A(n2965), .Z(n2972) );
  BUF_X1 U71 ( .A(n2920), .Z(n2925) );
  BUF_X1 U72 ( .A(n2965), .Z(n2971) );
  BUF_X1 U73 ( .A(n2921), .Z(n2926) );
  BUF_X1 U74 ( .A(n2921), .Z(n2927) );
  BUF_X1 U75 ( .A(n2921), .Z(n2928) );
  BUF_X1 U76 ( .A(n2964), .Z(n2968) );
  BUF_X1 U77 ( .A(n2965), .Z(n2970) );
  BUF_X1 U78 ( .A(n2964), .Z(n2969) );
  BUF_X1 U79 ( .A(n2966), .Z(n2974) );
  BUF_X1 U80 ( .A(n2966), .Z(n2973) );
  BUF_X1 U81 ( .A(n2922), .Z(n2930) );
  BUF_X1 U82 ( .A(n2922), .Z(n2929) );
  BUF_X1 U83 ( .A(n2838), .Z(n2845) );
  BUF_X1 U84 ( .A(n2838), .Z(n2844) );
  BUF_X1 U85 ( .A(n2838), .Z(n2843) );
  BUF_X1 U86 ( .A(n2975), .Z(n2978) );
  BUF_X1 U87 ( .A(n2839), .Z(n2847) );
  BUF_X1 U88 ( .A(n2839), .Z(n2846) );
  BUF_X1 U89 ( .A(n2953), .Z(n2957) );
  BUF_X1 U90 ( .A(n2953), .Z(n2956) );
  BUF_X1 U91 ( .A(n2976), .Z(n2983) );
  BUF_X1 U92 ( .A(n2976), .Z(n2982) );
  BUF_X1 U93 ( .A(n2975), .Z(n2979) );
  BUF_X1 U94 ( .A(n2976), .Z(n2981) );
  BUF_X1 U95 ( .A(n2975), .Z(n2980) );
  BUF_X1 U96 ( .A(n2977), .Z(n2985) );
  BUF_X1 U97 ( .A(n2977), .Z(n2984) );
  BUF_X1 U98 ( .A(n692), .Z(n3029) );
  BUF_X1 U99 ( .A(n694), .Z(n3023) );
  BUF_X1 U100 ( .A(n3008), .Z(n3011) );
  BUF_X1 U101 ( .A(n693), .Z(n3026) );
  BUF_X1 U102 ( .A(n2953), .Z(n2958) );
  BUF_X1 U103 ( .A(n2954), .Z(n2959) );
  BUF_X1 U104 ( .A(n2954), .Z(n2960) );
  BUF_X1 U105 ( .A(n2954), .Z(n2961) );
  BUF_X1 U106 ( .A(n2955), .Z(n2963) );
  BUF_X1 U107 ( .A(n2955), .Z(n2962) );
  BUF_X1 U108 ( .A(n1934), .Z(n2813) );
  BUF_X1 U109 ( .A(n1945), .Z(n2804) );
  BUF_X1 U110 ( .A(n1946), .Z(n2801) );
  BUF_X1 U111 ( .A(n2861), .Z(n2869) );
  BUF_X1 U112 ( .A(n1884), .Z(n2917) );
  BUF_X1 U113 ( .A(n681), .Z(n3039) );
  BUF_X1 U114 ( .A(n681), .Z(n3040) );
  BUF_X1 U115 ( .A(n681), .Z(n3041) );
  NAND2_X1 U116 ( .A1(n1867), .A2(read_address_2[0]), .ZN(n683) );
  BUF_X1 U117 ( .A(n696), .Z(n3015) );
  BUF_X1 U118 ( .A(n696), .Z(n3016) );
  NOR2_X1 U119 ( .A1(n2978), .A2(read_address_2[0]), .ZN(n693) );
  NOR2_X1 U120 ( .A1(n2967), .A2(read_address_2[0]), .ZN(n692) );
  NOR2_X1 U121 ( .A1(n1855), .A2(read_address_2[0]), .ZN(n694) );
  BUF_X1 U122 ( .A(n695), .Z(n3018) );
  BUF_X1 U123 ( .A(n697), .Z(n3012) );
  BUF_X1 U124 ( .A(n695), .Z(n3019) );
  BUF_X1 U125 ( .A(n697), .Z(n3013) );
  BUF_X1 U126 ( .A(n2892), .Z(n2895) );
  BUF_X1 U127 ( .A(n2892), .Z(n2896) );
  BUF_X1 U128 ( .A(n1884), .Z(n2918) );
  BUF_X1 U129 ( .A(n2892), .Z(n2897) );
  BUF_X1 U130 ( .A(n2893), .Z(n2900) );
  BUF_X1 U131 ( .A(n2893), .Z(n2899) );
  BUF_X1 U132 ( .A(n2893), .Z(n2898) );
  BUF_X1 U133 ( .A(n2894), .Z(n2902) );
  BUF_X1 U134 ( .A(n2894), .Z(n2901) );
  BUF_X1 U135 ( .A(n1932), .Z(n2814) );
  BUF_X1 U136 ( .A(n1943), .Z(n2805) );
  BUF_X1 U137 ( .A(n1932), .Z(n2815) );
  BUF_X1 U138 ( .A(n1943), .Z(n2806) );
  BUF_X1 U139 ( .A(n2881), .Z(n2884) );
  BUF_X1 U140 ( .A(n2881), .Z(n2885) );
  BUF_X1 U141 ( .A(n2881), .Z(n2886) );
  BUF_X1 U142 ( .A(n1910), .Z(n2914) );
  BUF_X1 U143 ( .A(n1923), .Z(n2823) );
  BUF_X1 U144 ( .A(n1910), .Z(n2915) );
  BUF_X1 U145 ( .A(n1923), .Z(n2824) );
  BUF_X1 U146 ( .A(n2882), .Z(n2889) );
  BUF_X1 U147 ( .A(n2882), .Z(n2888) );
  BUF_X1 U148 ( .A(n2882), .Z(n2887) );
  BUF_X1 U149 ( .A(n2931), .Z(n2934) );
  BUF_X1 U150 ( .A(n2826), .Z(n2829) );
  BUF_X1 U151 ( .A(n2870), .Z(n2873) );
  BUF_X1 U152 ( .A(n2826), .Z(n2830) );
  BUF_X1 U153 ( .A(n2870), .Z(n2874) );
  BUF_X1 U154 ( .A(n2883), .Z(n2891) );
  BUF_X1 U155 ( .A(n2883), .Z(n2890) );
  BUF_X1 U156 ( .A(n2932), .Z(n2939) );
  BUF_X1 U157 ( .A(n2932), .Z(n2938) );
  BUF_X1 U158 ( .A(n2931), .Z(n2935) );
  BUF_X1 U159 ( .A(n2932), .Z(n2937) );
  BUF_X1 U160 ( .A(n2931), .Z(n2936) );
  BUF_X1 U161 ( .A(n2933), .Z(n2941) );
  BUF_X1 U162 ( .A(n2933), .Z(n2940) );
  BUF_X1 U163 ( .A(n696), .Z(n3017) );
  BUF_X1 U164 ( .A(n1930), .Z(n2817) );
  BUF_X1 U165 ( .A(n1941), .Z(n2808) );
  BUF_X1 U166 ( .A(n1930), .Z(n2818) );
  BUF_X1 U167 ( .A(n1941), .Z(n2809) );
  BUF_X1 U168 ( .A(n2870), .Z(n2875) );
  BUF_X1 U169 ( .A(n2826), .Z(n2831) );
  BUF_X1 U170 ( .A(n695), .Z(n3020) );
  BUF_X1 U171 ( .A(n697), .Z(n3014) );
  BUF_X1 U172 ( .A(n2871), .Z(n2878) );
  BUF_X1 U173 ( .A(n2827), .Z(n2834) );
  BUF_X1 U174 ( .A(n2871), .Z(n2877) );
  BUF_X1 U175 ( .A(n2827), .Z(n2833) );
  BUF_X1 U176 ( .A(n2871), .Z(n2876) );
  BUF_X1 U177 ( .A(n2827), .Z(n2832) );
  BUF_X1 U178 ( .A(n2872), .Z(n2880) );
  BUF_X1 U179 ( .A(n2828), .Z(n2836) );
  BUF_X1 U180 ( .A(n2872), .Z(n2879) );
  BUF_X1 U181 ( .A(n2828), .Z(n2835) );
  BUF_X1 U182 ( .A(n1932), .Z(n2816) );
  BUF_X1 U183 ( .A(n1943), .Z(n2807) );
  BUF_X1 U184 ( .A(n1910), .Z(n2916) );
  BUF_X1 U185 ( .A(n1923), .Z(n2825) );
  BUF_X1 U186 ( .A(n1930), .Z(n2819) );
  BUF_X1 U187 ( .A(n1941), .Z(n2810) );
  BUF_X1 U188 ( .A(n1884), .Z(n2919) );
  NOR2_X1 U189 ( .A1(n2897), .A2(read_address_1[0]), .ZN(n1934) );
  NOR2_X1 U190 ( .A1(n2853), .A2(read_address_1[0]), .ZN(n1946) );
  NOR2_X1 U191 ( .A1(n2864), .A2(read_address_1[0]), .ZN(n1945) );
  BUF_X1 U192 ( .A(n698), .Z(n3008) );
  NOR2_X1 U193 ( .A1(n2934), .A2(read_address_2[0]), .ZN(n698) );
  INV_X1 U194 ( .A(n1855), .ZN(n702) );
  BUF_X1 U195 ( .A(n3042), .Z(n3046) );
  BUF_X1 U196 ( .A(n3042), .Z(n3044) );
  BUF_X1 U197 ( .A(n3042), .Z(n3045) );
  BUF_X1 U198 ( .A(n3043), .Z(n3047) );
  BUF_X1 U199 ( .A(n2369), .Z(n3050) );
  BUF_X1 U200 ( .A(n2369), .Z(n3049) );
  BUF_X1 U201 ( .A(n2365), .Z(n3053) );
  BUF_X1 U202 ( .A(n2365), .Z(n3052) );
  BUF_X1 U203 ( .A(n2361), .Z(n3056) );
  BUF_X1 U204 ( .A(n2361), .Z(n3055) );
  BUF_X1 U205 ( .A(n2357), .Z(n3059) );
  BUF_X1 U206 ( .A(n2357), .Z(n3058) );
  BUF_X1 U207 ( .A(n2353), .Z(n3062) );
  BUF_X1 U208 ( .A(n2353), .Z(n3061) );
  BUF_X1 U209 ( .A(n2349), .Z(n3065) );
  BUF_X1 U210 ( .A(n2349), .Z(n3064) );
  BUF_X1 U211 ( .A(n2345), .Z(n3068) );
  BUF_X1 U212 ( .A(n2345), .Z(n3067) );
  BUF_X1 U213 ( .A(n2341), .Z(n3071) );
  BUF_X1 U214 ( .A(n2341), .Z(n3070) );
  BUF_X1 U215 ( .A(n2337), .Z(n3074) );
  BUF_X1 U216 ( .A(n2337), .Z(n3073) );
  BUF_X1 U217 ( .A(n2333), .Z(n3077) );
  BUF_X1 U218 ( .A(n2333), .Z(n3076) );
  BUF_X1 U219 ( .A(n2329), .Z(n3080) );
  BUF_X1 U220 ( .A(n2329), .Z(n3079) );
  BUF_X1 U221 ( .A(n2325), .Z(n3083) );
  BUF_X1 U222 ( .A(n2325), .Z(n3082) );
  BUF_X1 U223 ( .A(n2321), .Z(n3086) );
  BUF_X1 U224 ( .A(n2321), .Z(n3085) );
  BUF_X1 U225 ( .A(n2317), .Z(n3089) );
  BUF_X1 U226 ( .A(n2317), .Z(n3088) );
  BUF_X1 U227 ( .A(n2313), .Z(n3092) );
  BUF_X1 U228 ( .A(n2313), .Z(n3091) );
  BUF_X1 U229 ( .A(n2309), .Z(n3095) );
  BUF_X1 U230 ( .A(n2309), .Z(n3094) );
  BUF_X1 U231 ( .A(n2305), .Z(n3098) );
  BUF_X1 U232 ( .A(n2305), .Z(n3097) );
  BUF_X1 U233 ( .A(n2301), .Z(n3101) );
  BUF_X1 U234 ( .A(n2301), .Z(n3100) );
  BUF_X1 U235 ( .A(n2297), .Z(n3104) );
  BUF_X1 U236 ( .A(n2297), .Z(n3103) );
  BUF_X1 U237 ( .A(n2293), .Z(n3107) );
  BUF_X1 U238 ( .A(n2293), .Z(n3106) );
  BUF_X1 U239 ( .A(n2289), .Z(n3110) );
  BUF_X1 U240 ( .A(n2289), .Z(n3109) );
  BUF_X1 U241 ( .A(n2285), .Z(n3113) );
  BUF_X1 U242 ( .A(n2285), .Z(n3112) );
  BUF_X1 U243 ( .A(n2281), .Z(n3116) );
  BUF_X1 U244 ( .A(n2281), .Z(n3115) );
  BUF_X1 U245 ( .A(n2277), .Z(n3119) );
  BUF_X1 U246 ( .A(n2277), .Z(n3118) );
  BUF_X1 U247 ( .A(n2273), .Z(n3122) );
  BUF_X1 U248 ( .A(n2273), .Z(n3121) );
  BUF_X1 U249 ( .A(n2269), .Z(n3125) );
  BUF_X1 U250 ( .A(n2269), .Z(n3124) );
  BUF_X1 U251 ( .A(n2265), .Z(n3128) );
  BUF_X1 U252 ( .A(n2265), .Z(n3127) );
  BUF_X1 U253 ( .A(n2261), .Z(n3131) );
  BUF_X1 U254 ( .A(n2261), .Z(n3130) );
  BUF_X1 U255 ( .A(n2257), .Z(n3134) );
  BUF_X1 U256 ( .A(n2257), .Z(n3133) );
  BUF_X1 U257 ( .A(n2253), .Z(n3137) );
  BUF_X1 U258 ( .A(n2253), .Z(n3136) );
  BUF_X1 U259 ( .A(n2249), .Z(n3140) );
  BUF_X1 U260 ( .A(n2249), .Z(n3139) );
  BUF_X1 U261 ( .A(n2369), .Z(n3051) );
  BUF_X1 U262 ( .A(n2365), .Z(n3054) );
  BUF_X1 U263 ( .A(n2361), .Z(n3057) );
  BUF_X1 U264 ( .A(n2357), .Z(n3060) );
  BUF_X1 U265 ( .A(n2353), .Z(n3063) );
  BUF_X1 U266 ( .A(n2349), .Z(n3066) );
  BUF_X1 U267 ( .A(n2345), .Z(n3069) );
  BUF_X1 U268 ( .A(n2341), .Z(n3072) );
  BUF_X1 U269 ( .A(n2337), .Z(n3075) );
  BUF_X1 U270 ( .A(n2333), .Z(n3078) );
  BUF_X1 U271 ( .A(n2329), .Z(n3081) );
  BUF_X1 U272 ( .A(n2325), .Z(n3084) );
  BUF_X1 U273 ( .A(n2321), .Z(n3087) );
  BUF_X1 U274 ( .A(n2317), .Z(n3090) );
  BUF_X1 U275 ( .A(n2313), .Z(n3093) );
  BUF_X1 U276 ( .A(n2309), .Z(n3096) );
  BUF_X1 U277 ( .A(n2305), .Z(n3099) );
  BUF_X1 U278 ( .A(n2301), .Z(n3102) );
  BUF_X1 U279 ( .A(n2297), .Z(n3105) );
  BUF_X1 U280 ( .A(n2293), .Z(n3108) );
  BUF_X1 U281 ( .A(n2289), .Z(n3111) );
  BUF_X1 U282 ( .A(n2285), .Z(n3114) );
  BUF_X1 U283 ( .A(n2281), .Z(n3117) );
  BUF_X1 U284 ( .A(n2277), .Z(n3120) );
  BUF_X1 U285 ( .A(n2273), .Z(n3123) );
  BUF_X1 U286 ( .A(n2269), .Z(n3126) );
  BUF_X1 U287 ( .A(n2265), .Z(n3129) );
  BUF_X1 U288 ( .A(n2261), .Z(n3132) );
  BUF_X1 U289 ( .A(n2257), .Z(n3135) );
  BUF_X1 U290 ( .A(n2253), .Z(n3138) );
  BUF_X1 U291 ( .A(n2249), .Z(n3141) );
  BUF_X1 U292 ( .A(n3043), .Z(n3048) );
  INV_X1 U293 ( .A(n3241), .ZN(n3240) );
  BUF_X1 U294 ( .A(n685), .Z(n3033) );
  BUF_X1 U295 ( .A(n685), .Z(n3034) );
  BUF_X1 U296 ( .A(n687), .Z(n3030) );
  BUF_X1 U297 ( .A(n685), .Z(n3035) );
  NOR2_X1 U298 ( .A1(n1879), .A2(n3030), .ZN(n1867) );
  NAND2_X1 U299 ( .A1(n1867), .A2(n3239), .ZN(n681) );
  INV_X1 U300 ( .A(n2772), .ZN(n1884) );
  OAI221_X1 U301 ( .B1(n921), .B2(n3041), .C1(n922), .C2(n3038), .A(n923), 
        .ZN(data_reg_2[3]) );
  NOR4_X1 U302 ( .A1(n938), .A2(n939), .A3(n940), .A4(n941), .ZN(n922) );
  NOR4_X1 U303 ( .A1(n948), .A2(n949), .A3(n950), .A4(n951), .ZN(n921) );
  OAI221_X1 U304 ( .B1(n884), .B2(n3041), .C1(n885), .C2(n3038), .A(n886), 
        .ZN(data_reg_2[4]) );
  NOR4_X1 U305 ( .A1(n901), .A2(n902), .A3(n903), .A4(n904), .ZN(n885) );
  NOR4_X1 U306 ( .A1(n911), .A2(n912), .A3(n913), .A4(n914), .ZN(n884) );
  OAI221_X1 U307 ( .B1(n847), .B2(n3041), .C1(n848), .C2(n3038), .A(n849), 
        .ZN(data_reg_2[5]) );
  NOR4_X1 U308 ( .A1(n864), .A2(n865), .A3(n866), .A4(n867), .ZN(n848) );
  NOR4_X1 U309 ( .A1(n874), .A2(n875), .A3(n876), .A4(n877), .ZN(n847) );
  OAI221_X1 U310 ( .B1(n810), .B2(n3041), .C1(n811), .C2(n3038), .A(n812), 
        .ZN(data_reg_2[6]) );
  NOR4_X1 U311 ( .A1(n827), .A2(n828), .A3(n829), .A4(n830), .ZN(n811) );
  NOR4_X1 U312 ( .A1(n837), .A2(n838), .A3(n839), .A4(n840), .ZN(n810) );
  OAI221_X1 U313 ( .B1(n773), .B2(n3041), .C1(n774), .C2(n3038), .A(n775), 
        .ZN(data_reg_2[7]) );
  NOR4_X1 U314 ( .A1(n800), .A2(n801), .A3(n802), .A4(n803), .ZN(n773) );
  NOR4_X1 U315 ( .A1(n790), .A2(n791), .A3(n792), .A4(n793), .ZN(n774) );
  OAI221_X1 U316 ( .B1(n736), .B2(n3041), .C1(n737), .C2(n3038), .A(n738), 
        .ZN(data_reg_2[8]) );
  NOR4_X1 U317 ( .A1(n753), .A2(n754), .A3(n755), .A4(n756), .ZN(n737) );
  NOR4_X1 U318 ( .A1(n763), .A2(n764), .A3(n765), .A4(n766), .ZN(n736) );
  OAI221_X1 U319 ( .B1(n680), .B2(n3041), .C1(n682), .C2(n3038), .A(n684), 
        .ZN(data_reg_2[9]) );
  NOR4_X1 U320 ( .A1(n716), .A2(n717), .A3(n718), .A4(n719), .ZN(n682) );
  NOR4_X1 U321 ( .A1(n726), .A2(n727), .A3(n728), .A4(n729), .ZN(n680) );
  OAI221_X1 U322 ( .B1(n958), .B2(n3041), .C1(n959), .C2(n3038), .A(n960), 
        .ZN(data_reg_2[31]) );
  NOR4_X1 U323 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .ZN(n959) );
  NOR4_X1 U324 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n958) );
  OAI221_X1 U325 ( .B1(n1846), .B2(n3039), .C1(n1847), .C2(n3036), .A(n1848), 
        .ZN(data_reg_2[0]) );
  NOR4_X1 U326 ( .A1(n1868), .A2(n1869), .A3(n1870), .A4(n1871), .ZN(n1847) );
  NOR4_X1 U327 ( .A1(n1889), .A2(n1890), .A3(n1891), .A4(n1892), .ZN(n1846) );
  OAI221_X1 U328 ( .B1(n1439), .B2(n3039), .C1(n1440), .C2(n3036), .A(n1441), 
        .ZN(data_reg_2[1]) );
  NOR4_X1 U329 ( .A1(n1456), .A2(n1457), .A3(n1458), .A4(n1459), .ZN(n1440) );
  NOR4_X1 U330 ( .A1(n1466), .A2(n1467), .A3(n1468), .A4(n1469), .ZN(n1439) );
  OAI221_X1 U331 ( .B1(n1032), .B2(n3040), .C1(n1033), .C2(n3037), .A(n1034), 
        .ZN(data_reg_2[2]) );
  NOR4_X1 U332 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1033) );
  NOR4_X1 U333 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1032) );
  OAI221_X1 U334 ( .B1(n1809), .B2(n3039), .C1(n1810), .C2(n3036), .A(n1811), 
        .ZN(data_reg_2[10]) );
  NOR4_X1 U335 ( .A1(n1836), .A2(n1837), .A3(n1838), .A4(n1839), .ZN(n1809) );
  NOR4_X1 U336 ( .A1(n1826), .A2(n1827), .A3(n1828), .A4(n1829), .ZN(n1810) );
  OAI221_X1 U337 ( .B1(n1772), .B2(n3039), .C1(n1773), .C2(n3036), .A(n1774), 
        .ZN(data_reg_2[11]) );
  NOR4_X1 U338 ( .A1(n1789), .A2(n1790), .A3(n1791), .A4(n1792), .ZN(n1773) );
  NOR4_X1 U339 ( .A1(n1799), .A2(n1800), .A3(n1801), .A4(n1802), .ZN(n1772) );
  OAI221_X1 U340 ( .B1(n1735), .B2(n3039), .C1(n1736), .C2(n3036), .A(n1737), 
        .ZN(data_reg_2[12]) );
  NOR4_X1 U341 ( .A1(n1752), .A2(n1753), .A3(n1754), .A4(n1755), .ZN(n1736) );
  NOR4_X1 U342 ( .A1(n1762), .A2(n1763), .A3(n1764), .A4(n1765), .ZN(n1735) );
  OAI221_X1 U343 ( .B1(n1698), .B2(n3039), .C1(n1699), .C2(n3036), .A(n1700), 
        .ZN(data_reg_2[13]) );
  NOR4_X1 U344 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(n1698) );
  NOR4_X1 U345 ( .A1(n1715), .A2(n1716), .A3(n1717), .A4(n1718), .ZN(n1699) );
  OAI221_X1 U346 ( .B1(n1661), .B2(n3039), .C1(n1662), .C2(n3036), .A(n1663), 
        .ZN(data_reg_2[14]) );
  NOR4_X1 U347 ( .A1(n1678), .A2(n1679), .A3(n1680), .A4(n1681), .ZN(n1662) );
  NOR4_X1 U348 ( .A1(n1688), .A2(n1689), .A3(n1690), .A4(n1691), .ZN(n1661) );
  OAI221_X1 U349 ( .B1(n1624), .B2(n3039), .C1(n1625), .C2(n3036), .A(n1626), 
        .ZN(data_reg_2[15]) );
  NOR4_X1 U350 ( .A1(n1641), .A2(n1642), .A3(n1643), .A4(n1644), .ZN(n1625) );
  NOR4_X1 U351 ( .A1(n1651), .A2(n1652), .A3(n1653), .A4(n1654), .ZN(n1624) );
  OAI221_X1 U352 ( .B1(n1587), .B2(n3039), .C1(n1588), .C2(n3036), .A(n1589), 
        .ZN(data_reg_2[16]) );
  NOR4_X1 U353 ( .A1(n1604), .A2(n1605), .A3(n1606), .A4(n1607), .ZN(n1588) );
  NOR4_X1 U354 ( .A1(n1614), .A2(n1615), .A3(n1616), .A4(n1617), .ZN(n1587) );
  OAI221_X1 U355 ( .B1(n1550), .B2(n3039), .C1(n1551), .C2(n3036), .A(n1552), 
        .ZN(data_reg_2[17]) );
  NOR4_X1 U356 ( .A1(n1567), .A2(n1568), .A3(n1569), .A4(n1570), .ZN(n1551) );
  NOR4_X1 U357 ( .A1(n1577), .A2(n1578), .A3(n1579), .A4(n1580), .ZN(n1550) );
  OAI221_X1 U358 ( .B1(n1513), .B2(n3039), .C1(n1514), .C2(n3036), .A(n1515), 
        .ZN(data_reg_2[18]) );
  NOR4_X1 U359 ( .A1(n1530), .A2(n1531), .A3(n1532), .A4(n1533), .ZN(n1514) );
  NOR4_X1 U360 ( .A1(n1540), .A2(n1541), .A3(n1542), .A4(n1543), .ZN(n1513) );
  OAI221_X1 U361 ( .B1(n1476), .B2(n3039), .C1(n1477), .C2(n3036), .A(n1478), 
        .ZN(data_reg_2[19]) );
  NOR4_X1 U362 ( .A1(n1493), .A2(n1494), .A3(n1495), .A4(n1496), .ZN(n1477) );
  NOR4_X1 U363 ( .A1(n1503), .A2(n1504), .A3(n1505), .A4(n1506), .ZN(n1476) );
  OAI221_X1 U364 ( .B1(n1402), .B2(n3040), .C1(n1403), .C2(n3037), .A(n1404), 
        .ZN(data_reg_2[20]) );
  NOR4_X1 U365 ( .A1(n1419), .A2(n1420), .A3(n1421), .A4(n1422), .ZN(n1403) );
  NOR4_X1 U366 ( .A1(n1429), .A2(n1430), .A3(n1431), .A4(n1432), .ZN(n1402) );
  OAI221_X1 U367 ( .B1(n1365), .B2(n3040), .C1(n1366), .C2(n3037), .A(n1367), 
        .ZN(data_reg_2[21]) );
  NOR4_X1 U368 ( .A1(n1382), .A2(n1383), .A3(n1384), .A4(n1385), .ZN(n1366) );
  NOR4_X1 U369 ( .A1(n1392), .A2(n1393), .A3(n1394), .A4(n1395), .ZN(n1365) );
  OAI221_X1 U370 ( .B1(n1328), .B2(n3040), .C1(n1329), .C2(n3037), .A(n1330), 
        .ZN(data_reg_2[22]) );
  NOR4_X1 U371 ( .A1(n1345), .A2(n1346), .A3(n1347), .A4(n1348), .ZN(n1329) );
  NOR4_X1 U372 ( .A1(n1355), .A2(n1356), .A3(n1357), .A4(n1358), .ZN(n1328) );
  OAI221_X1 U373 ( .B1(n1291), .B2(n3040), .C1(n1292), .C2(n3037), .A(n1293), 
        .ZN(data_reg_2[23]) );
  NOR4_X1 U374 ( .A1(n1308), .A2(n1309), .A3(n1310), .A4(n1311), .ZN(n1292) );
  NOR4_X1 U375 ( .A1(n1318), .A2(n1319), .A3(n1320), .A4(n1321), .ZN(n1291) );
  OAI221_X1 U376 ( .B1(n1254), .B2(n3040), .C1(n1255), .C2(n3037), .A(n1256), 
        .ZN(data_reg_2[24]) );
  NOR4_X1 U377 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1255) );
  NOR4_X1 U378 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1254) );
  OAI221_X1 U379 ( .B1(n1217), .B2(n3040), .C1(n1218), .C2(n3037), .A(n1219), 
        .ZN(data_reg_2[25]) );
  NOR4_X1 U380 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1218) );
  NOR4_X1 U381 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1217) );
  OAI221_X1 U382 ( .B1(n1180), .B2(n3040), .C1(n1181), .C2(n3037), .A(n1182), 
        .ZN(data_reg_2[26]) );
  NOR4_X1 U383 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1181) );
  NOR4_X1 U384 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1180) );
  OAI221_X1 U385 ( .B1(n1143), .B2(n3040), .C1(n1144), .C2(n3037), .A(n1145), 
        .ZN(data_reg_2[27]) );
  NOR4_X1 U386 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1144) );
  NOR4_X1 U387 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1143) );
  OAI221_X1 U388 ( .B1(n1106), .B2(n3040), .C1(n1107), .C2(n3037), .A(n1108), 
        .ZN(data_reg_2[28]) );
  NOR4_X1 U389 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1107) );
  NOR4_X1 U390 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1106) );
  OAI221_X1 U391 ( .B1(n1069), .B2(n3040), .C1(n1070), .C2(n3037), .A(n1071), 
        .ZN(data_reg_2[29]) );
  NOR4_X1 U392 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1070) );
  NOR4_X1 U393 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1069) );
  OAI221_X1 U394 ( .B1(n995), .B2(n3040), .C1(n996), .C2(n3037), .A(n997), 
        .ZN(data_reg_2[30]) );
  NOR4_X1 U395 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n996) );
  NOR4_X1 U396 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n995) );
  INV_X1 U397 ( .A(n3239), .ZN(n3238) );
  BUF_X1 U398 ( .A(n1928), .Z(n2820) );
  BUF_X1 U399 ( .A(n1928), .Z(n2821) );
  OAI22_X1 U400 ( .A1(n2934), .A2(n1893), .B1(n2923), .B2(n1894), .ZN(n1892)
         );
  OAI22_X1 U401 ( .A1(n2933), .A2(n1872), .B1(n2923), .B2(n1873), .ZN(n1871)
         );
  OAI22_X1 U402 ( .A1(n2939), .A2(n1470), .B1(n2925), .B2(n1471), .ZN(n1469)
         );
  OAI22_X1 U403 ( .A1(n2939), .A2(n1460), .B1(n2925), .B2(n1461), .ZN(n1459)
         );
  OAI22_X1 U404 ( .A1(n2936), .A2(n1063), .B1(n2928), .B2(n1064), .ZN(n1062)
         );
  OAI22_X1 U405 ( .A1(n2936), .A2(n1053), .B1(n2928), .B2(n1054), .ZN(n1052)
         );
  OAI22_X1 U406 ( .A1(n2935), .A2(n952), .B1(n2929), .B2(n953), .ZN(n951) );
  OAI22_X1 U407 ( .A1(n2935), .A2(n942), .B1(n2929), .B2(n943), .ZN(n941) );
  OAI22_X1 U408 ( .A1(n2935), .A2(n915), .B1(n2929), .B2(n916), .ZN(n914) );
  OAI22_X1 U409 ( .A1(n2935), .A2(n905), .B1(n2929), .B2(n906), .ZN(n904) );
  OAI22_X1 U410 ( .A1(n2935), .A2(n878), .B1(n2929), .B2(n879), .ZN(n877) );
  OAI22_X1 U411 ( .A1(n2935), .A2(n868), .B1(n2929), .B2(n869), .ZN(n867) );
  OAI22_X1 U412 ( .A1(n2935), .A2(n841), .B1(n2930), .B2(n842), .ZN(n840) );
  OAI22_X1 U413 ( .A1(n2934), .A2(n831), .B1(n2930), .B2(n832), .ZN(n830) );
  OAI22_X1 U414 ( .A1(n2934), .A2(n794), .B1(n2930), .B2(n795), .ZN(n793) );
  OAI22_X1 U415 ( .A1(n2934), .A2(n804), .B1(n2930), .B2(n805), .ZN(n803) );
  OAI22_X1 U416 ( .A1(n2934), .A2(n767), .B1(n2930), .B2(n768), .ZN(n766) );
  OAI22_X1 U417 ( .A1(n2934), .A2(n757), .B1(n2930), .B2(n758), .ZN(n756) );
  OAI22_X1 U418 ( .A1(n2934), .A2(n730), .B1(n2930), .B2(n731), .ZN(n729) );
  OAI22_X1 U419 ( .A1(n2934), .A2(n720), .B1(n2930), .B2(n721), .ZN(n719) );
  OAI22_X1 U420 ( .A1(n2941), .A2(n1830), .B1(n2923), .B2(n1831), .ZN(n1829)
         );
  OAI22_X1 U421 ( .A1(n2941), .A2(n1840), .B1(n2923), .B2(n1841), .ZN(n1839)
         );
  OAI22_X1 U422 ( .A1(n2941), .A2(n1803), .B1(n2923), .B2(n1804), .ZN(n1802)
         );
  OAI22_X1 U423 ( .A1(n2941), .A2(n1793), .B1(n2923), .B2(n1794), .ZN(n1792)
         );
  OAI22_X1 U424 ( .A1(n2941), .A2(n1766), .B1(n2923), .B2(n1767), .ZN(n1765)
         );
  OAI22_X1 U425 ( .A1(n2941), .A2(n1756), .B1(n2923), .B2(n1757), .ZN(n1755)
         );
  OAI22_X1 U426 ( .A1(n2941), .A2(n1719), .B1(n2924), .B2(n1720), .ZN(n1718)
         );
  OAI22_X1 U427 ( .A1(n2941), .A2(n1729), .B1(n2924), .B2(n1730), .ZN(n1728)
         );
  OAI22_X1 U428 ( .A1(n2940), .A2(n1692), .B1(n2924), .B2(n1693), .ZN(n1691)
         );
  OAI22_X1 U429 ( .A1(n2940), .A2(n1682), .B1(n2924), .B2(n1683), .ZN(n1681)
         );
  OAI22_X1 U430 ( .A1(n2940), .A2(n1655), .B1(n2924), .B2(n1656), .ZN(n1654)
         );
  OAI22_X1 U431 ( .A1(n2940), .A2(n1645), .B1(n2924), .B2(n1646), .ZN(n1644)
         );
  OAI22_X1 U432 ( .A1(n2940), .A2(n1618), .B1(n2924), .B2(n1619), .ZN(n1617)
         );
  OAI22_X1 U433 ( .A1(n2940), .A2(n1608), .B1(n2924), .B2(n1609), .ZN(n1607)
         );
  OAI22_X1 U434 ( .A1(n2940), .A2(n1581), .B1(n2925), .B2(n1582), .ZN(n1580)
         );
  OAI22_X1 U435 ( .A1(n2940), .A2(n1571), .B1(n2925), .B2(n1572), .ZN(n1570)
         );
  OAI22_X1 U436 ( .A1(n2939), .A2(n1544), .B1(n2925), .B2(n1545), .ZN(n1543)
         );
  OAI22_X1 U437 ( .A1(n2939), .A2(n1534), .B1(n2925), .B2(n1535), .ZN(n1533)
         );
  OAI22_X1 U438 ( .A1(n2939), .A2(n1507), .B1(n2925), .B2(n1508), .ZN(n1506)
         );
  OAI22_X1 U439 ( .A1(n2939), .A2(n1497), .B1(n2925), .B2(n1498), .ZN(n1496)
         );
  OAI22_X1 U440 ( .A1(n2939), .A2(n1433), .B1(n2926), .B2(n1434), .ZN(n1432)
         );
  OAI22_X1 U441 ( .A1(n2939), .A2(n1423), .B1(n2926), .B2(n1424), .ZN(n1422)
         );
  OAI22_X1 U442 ( .A1(n2938), .A2(n1396), .B1(n2926), .B2(n1397), .ZN(n1395)
         );
  OAI22_X1 U443 ( .A1(n2938), .A2(n1386), .B1(n2926), .B2(n1387), .ZN(n1385)
         );
  OAI22_X1 U444 ( .A1(n2938), .A2(n1359), .B1(n2926), .B2(n1360), .ZN(n1358)
         );
  OAI22_X1 U445 ( .A1(n2938), .A2(n1349), .B1(n2926), .B2(n1350), .ZN(n1348)
         );
  OAI22_X1 U446 ( .A1(n2938), .A2(n1322), .B1(n2926), .B2(n1323), .ZN(n1321)
         );
  OAI22_X1 U447 ( .A1(n2938), .A2(n1312), .B1(n2926), .B2(n1313), .ZN(n1311)
         );
  OAI22_X1 U448 ( .A1(n2938), .A2(n1285), .B1(n2927), .B2(n1286), .ZN(n1284)
         );
  OAI22_X1 U449 ( .A1(n2937), .A2(n1275), .B1(n2927), .B2(n1276), .ZN(n1274)
         );
  OAI22_X1 U450 ( .A1(n2937), .A2(n1248), .B1(n2927), .B2(n1249), .ZN(n1247)
         );
  OAI22_X1 U451 ( .A1(n2937), .A2(n1238), .B1(n2927), .B2(n1239), .ZN(n1237)
         );
  OAI22_X1 U452 ( .A1(n2937), .A2(n1211), .B1(n2927), .B2(n1212), .ZN(n1210)
         );
  OAI22_X1 U453 ( .A1(n2937), .A2(n1201), .B1(n2927), .B2(n1202), .ZN(n1200)
         );
  OAI22_X1 U454 ( .A1(n2937), .A2(n1174), .B1(n2927), .B2(n1175), .ZN(n1173)
         );
  OAI22_X1 U455 ( .A1(n2937), .A2(n1164), .B1(n2927), .B2(n1165), .ZN(n1163)
         );
  OAI22_X1 U456 ( .A1(n2937), .A2(n1137), .B1(n2928), .B2(n1138), .ZN(n1136)
         );
  OAI22_X1 U457 ( .A1(n2936), .A2(n1127), .B1(n2928), .B2(n1128), .ZN(n1126)
         );
  OAI22_X1 U458 ( .A1(n2936), .A2(n1100), .B1(n2928), .B2(n1101), .ZN(n1099)
         );
  OAI22_X1 U459 ( .A1(n2936), .A2(n1090), .B1(n2928), .B2(n1091), .ZN(n1089)
         );
  OAI22_X1 U460 ( .A1(n2936), .A2(n1026), .B1(n2928), .B2(n1027), .ZN(n1025)
         );
  OAI22_X1 U461 ( .A1(n2936), .A2(n1016), .B1(n2928), .B2(n1017), .ZN(n1015)
         );
  OAI22_X1 U462 ( .A1(n2936), .A2(n989), .B1(n2929), .B2(n990), .ZN(n988) );
  OAI22_X1 U463 ( .A1(n2935), .A2(n979), .B1(n2929), .B2(n980), .ZN(n978) );
  OAI22_X1 U464 ( .A1(n2985), .A2(n1862), .B1(n2974), .B2(n1863), .ZN(n1861)
         );
  OAI22_X1 U465 ( .A1(n2941), .A2(n1865), .B1(n2923), .B2(n1866), .ZN(n1864)
         );
  OAI22_X1 U466 ( .A1(n2983), .A2(n1451), .B1(n2972), .B2(n1452), .ZN(n1450)
         );
  OAI22_X1 U467 ( .A1(n2939), .A2(n1454), .B1(n2925), .B2(n1455), .ZN(n1453)
         );
  OAI22_X1 U468 ( .A1(n2980), .A2(n1044), .B1(n2969), .B2(n1045), .ZN(n1043)
         );
  OAI22_X1 U469 ( .A1(n2936), .A2(n1047), .B1(n2928), .B2(n1048), .ZN(n1046)
         );
  OAI22_X1 U470 ( .A1(n2979), .A2(n933), .B1(n2968), .B2(n934), .ZN(n932) );
  OAI22_X1 U471 ( .A1(n2935), .A2(n936), .B1(n2929), .B2(n937), .ZN(n935) );
  OAI22_X1 U472 ( .A1(n2979), .A2(n896), .B1(n2968), .B2(n897), .ZN(n895) );
  OAI22_X1 U473 ( .A1(n2935), .A2(n899), .B1(n2929), .B2(n900), .ZN(n898) );
  OAI22_X1 U474 ( .A1(n2979), .A2(n859), .B1(n2968), .B2(n860), .ZN(n858) );
  OAI22_X1 U475 ( .A1(n2935), .A2(n862), .B1(n2929), .B2(n863), .ZN(n861) );
  OAI22_X1 U476 ( .A1(n2978), .A2(n822), .B1(n2967), .B2(n823), .ZN(n821) );
  OAI22_X1 U477 ( .A1(n2934), .A2(n825), .B1(n2930), .B2(n826), .ZN(n824) );
  OAI22_X1 U478 ( .A1(n2978), .A2(n785), .B1(n2967), .B2(n786), .ZN(n784) );
  OAI22_X1 U479 ( .A1(n2934), .A2(n788), .B1(n2930), .B2(n789), .ZN(n787) );
  OAI22_X1 U480 ( .A1(n2978), .A2(n748), .B1(n2967), .B2(n749), .ZN(n747) );
  OAI22_X1 U481 ( .A1(n2934), .A2(n751), .B1(n2930), .B2(n752), .ZN(n750) );
  OAI22_X1 U482 ( .A1(n2982), .A2(n706), .B1(n2971), .B2(n708), .ZN(n704) );
  OAI22_X1 U483 ( .A1(n2938), .A2(n713), .B1(n2930), .B2(n715), .ZN(n711) );
  OAI22_X1 U484 ( .A1(n2985), .A2(n1821), .B1(n2974), .B2(n1822), .ZN(n1820)
         );
  OAI22_X1 U485 ( .A1(n2941), .A2(n1824), .B1(n2923), .B2(n1825), .ZN(n1823)
         );
  OAI22_X1 U486 ( .A1(n2985), .A2(n1784), .B1(n2974), .B2(n1785), .ZN(n1783)
         );
  OAI22_X1 U487 ( .A1(n2941), .A2(n1787), .B1(n2923), .B2(n1788), .ZN(n1786)
         );
  OAI22_X1 U488 ( .A1(n2985), .A2(n1747), .B1(n2974), .B2(n1748), .ZN(n1746)
         );
  OAI22_X1 U489 ( .A1(n2941), .A2(n1750), .B1(n2923), .B2(n1751), .ZN(n1749)
         );
  OAI22_X1 U490 ( .A1(n2984), .A2(n1710), .B1(n2973), .B2(n1711), .ZN(n1709)
         );
  OAI22_X1 U491 ( .A1(n2940), .A2(n1713), .B1(n2924), .B2(n1714), .ZN(n1712)
         );
  OAI22_X1 U492 ( .A1(n2984), .A2(n1673), .B1(n2973), .B2(n1674), .ZN(n1672)
         );
  OAI22_X1 U493 ( .A1(n2940), .A2(n1676), .B1(n2924), .B2(n1677), .ZN(n1675)
         );
  OAI22_X1 U494 ( .A1(n2984), .A2(n1636), .B1(n2973), .B2(n1637), .ZN(n1635)
         );
  OAI22_X1 U495 ( .A1(n2940), .A2(n1639), .B1(n2924), .B2(n1640), .ZN(n1638)
         );
  OAI22_X1 U496 ( .A1(n2984), .A2(n1599), .B1(n2973), .B2(n1600), .ZN(n1598)
         );
  OAI22_X1 U497 ( .A1(n2940), .A2(n1602), .B1(n2924), .B2(n1603), .ZN(n1601)
         );
  OAI22_X1 U498 ( .A1(n2983), .A2(n1562), .B1(n2972), .B2(n1563), .ZN(n1561)
         );
  OAI22_X1 U499 ( .A1(n2939), .A2(n1565), .B1(n2925), .B2(n1566), .ZN(n1564)
         );
  OAI22_X1 U500 ( .A1(n2983), .A2(n1525), .B1(n2972), .B2(n1526), .ZN(n1524)
         );
  OAI22_X1 U501 ( .A1(n2939), .A2(n1528), .B1(n2925), .B2(n1529), .ZN(n1527)
         );
  OAI22_X1 U502 ( .A1(n2983), .A2(n1488), .B1(n2972), .B2(n1489), .ZN(n1487)
         );
  OAI22_X1 U503 ( .A1(n2939), .A2(n1491), .B1(n2925), .B2(n1492), .ZN(n1490)
         );
  OAI22_X1 U504 ( .A1(n2982), .A2(n1414), .B1(n2971), .B2(n1415), .ZN(n1413)
         );
  OAI22_X1 U505 ( .A1(n2938), .A2(n1417), .B1(n2926), .B2(n1418), .ZN(n1416)
         );
  OAI22_X1 U506 ( .A1(n2982), .A2(n1377), .B1(n2971), .B2(n1378), .ZN(n1376)
         );
  OAI22_X1 U507 ( .A1(n2938), .A2(n1380), .B1(n2926), .B2(n1381), .ZN(n1379)
         );
  OAI22_X1 U508 ( .A1(n2982), .A2(n1340), .B1(n2971), .B2(n1341), .ZN(n1339)
         );
  OAI22_X1 U509 ( .A1(n2938), .A2(n1343), .B1(n2926), .B2(n1344), .ZN(n1342)
         );
  OAI22_X1 U510 ( .A1(n2982), .A2(n1303), .B1(n2971), .B2(n1304), .ZN(n1302)
         );
  OAI22_X1 U511 ( .A1(n2938), .A2(n1306), .B1(n2926), .B2(n1307), .ZN(n1305)
         );
  OAI22_X1 U512 ( .A1(n2981), .A2(n1266), .B1(n2970), .B2(n1267), .ZN(n1265)
         );
  OAI22_X1 U513 ( .A1(n2937), .A2(n1269), .B1(n2927), .B2(n1270), .ZN(n1268)
         );
  OAI22_X1 U514 ( .A1(n2981), .A2(n1229), .B1(n2970), .B2(n1230), .ZN(n1228)
         );
  OAI22_X1 U515 ( .A1(n2937), .A2(n1232), .B1(n2927), .B2(n1233), .ZN(n1231)
         );
  OAI22_X1 U516 ( .A1(n2981), .A2(n1192), .B1(n2970), .B2(n1193), .ZN(n1191)
         );
  OAI22_X1 U517 ( .A1(n2937), .A2(n1195), .B1(n2927), .B2(n1196), .ZN(n1194)
         );
  OAI22_X1 U518 ( .A1(n2981), .A2(n1155), .B1(n2970), .B2(n1156), .ZN(n1154)
         );
  OAI22_X1 U519 ( .A1(n2937), .A2(n1158), .B1(n2927), .B2(n1159), .ZN(n1157)
         );
  OAI22_X1 U520 ( .A1(n2980), .A2(n1118), .B1(n2969), .B2(n1119), .ZN(n1117)
         );
  OAI22_X1 U521 ( .A1(n2936), .A2(n1121), .B1(n2928), .B2(n1122), .ZN(n1120)
         );
  OAI22_X1 U522 ( .A1(n2980), .A2(n1081), .B1(n2969), .B2(n1082), .ZN(n1080)
         );
  OAI22_X1 U523 ( .A1(n2936), .A2(n1084), .B1(n2928), .B2(n1085), .ZN(n1083)
         );
  OAI22_X1 U524 ( .A1(n2980), .A2(n1007), .B1(n2969), .B2(n1008), .ZN(n1006)
         );
  OAI22_X1 U525 ( .A1(n2936), .A2(n1010), .B1(n2928), .B2(n1011), .ZN(n1009)
         );
  OAI22_X1 U526 ( .A1(n2979), .A2(n970), .B1(n2968), .B2(n971), .ZN(n969) );
  OAI22_X1 U527 ( .A1(n2935), .A2(n973), .B1(n2929), .B2(n974), .ZN(n972) );
  OAI22_X1 U528 ( .A1(n1862), .A2(n2851), .B1(n1863), .B2(n2862), .ZN(n2783)
         );
  OAI22_X1 U529 ( .A1(n1865), .A2(n2895), .B1(n1866), .B2(n2906), .ZN(n2784)
         );
  OAI22_X1 U530 ( .A1(n1451), .A2(n2852), .B1(n1452), .B2(n2863), .ZN(n2505)
         );
  OAI22_X1 U531 ( .A1(n1454), .A2(n2896), .B1(n1455), .B2(n2907), .ZN(n2506)
         );
  OAI22_X1 U532 ( .A1(n1044), .A2(n2853), .B1(n1045), .B2(n2864), .ZN(n2175)
         );
  OAI22_X1 U533 ( .A1(n1047), .A2(n2897), .B1(n1048), .B2(n2908), .ZN(n2177)
         );
  OAI22_X1 U534 ( .A1(n933), .A2(n2851), .B1(n934), .B2(n2862), .ZN(n2092) );
  OAI22_X1 U535 ( .A1(n936), .A2(n2895), .B1(n937), .B2(n2907), .ZN(n2093) );
  OAI22_X1 U536 ( .A1(n896), .A2(n2852), .B1(n897), .B2(n2863), .ZN(n2067) );
  OAI22_X1 U537 ( .A1(n899), .A2(n2896), .B1(n900), .B2(n2907), .ZN(n2068) );
  OAI22_X1 U538 ( .A1(n859), .A2(n2851), .B1(n860), .B2(n2862), .ZN(n2042) );
  OAI22_X1 U539 ( .A1(n862), .A2(n2895), .B1(n863), .B2(n2907), .ZN(n2043) );
  OAI22_X1 U540 ( .A1(n822), .A2(n2852), .B1(n823), .B2(n2863), .ZN(n2017) );
  OAI22_X1 U541 ( .A1(n825), .A2(n2896), .B1(n826), .B2(n2906), .ZN(n2018) );
  OAI22_X1 U542 ( .A1(n785), .A2(n2851), .B1(n786), .B2(n2862), .ZN(n1992) );
  OAI22_X1 U543 ( .A1(n788), .A2(n2895), .B1(n789), .B2(n2906), .ZN(n1993) );
  OAI22_X1 U544 ( .A1(n748), .A2(n2851), .B1(n749), .B2(n2862), .ZN(n1967) );
  OAI22_X1 U545 ( .A1(n751), .A2(n2895), .B1(n752), .B2(n2906), .ZN(n1968) );
  OAI22_X1 U546 ( .A1(n706), .A2(n2851), .B1(n708), .B2(n2862), .ZN(n1938) );
  OAI22_X1 U547 ( .A1(n713), .A2(n2895), .B1(n715), .B2(n2906), .ZN(n1939) );
  OAI22_X1 U548 ( .A1(n1821), .A2(n2851), .B1(n1822), .B2(n2862), .ZN(n2755)
         );
  OAI22_X1 U549 ( .A1(n1824), .A2(n2895), .B1(n1825), .B2(n2906), .ZN(n2756)
         );
  OAI22_X1 U550 ( .A1(n1784), .A2(n2851), .B1(n1785), .B2(n2862), .ZN(n2730)
         );
  OAI22_X1 U551 ( .A1(n1787), .A2(n2895), .B1(n1788), .B2(n2906), .ZN(n2731)
         );
  OAI22_X1 U552 ( .A1(n1747), .A2(n2851), .B1(n1748), .B2(n2862), .ZN(n2705)
         );
  OAI22_X1 U553 ( .A1(n1750), .A2(n2895), .B1(n1751), .B2(n2906), .ZN(n2706)
         );
  OAI22_X1 U554 ( .A1(n1710), .A2(n2851), .B1(n1711), .B2(n2862), .ZN(n2680)
         );
  OAI22_X1 U555 ( .A1(n1713), .A2(n2895), .B1(n1714), .B2(n2906), .ZN(n2681)
         );
  OAI22_X1 U556 ( .A1(n1673), .A2(n2851), .B1(n1674), .B2(n2862), .ZN(n2655)
         );
  OAI22_X1 U557 ( .A1(n1676), .A2(n2895), .B1(n1677), .B2(n2906), .ZN(n2656)
         );
  OAI22_X1 U558 ( .A1(n1636), .A2(n2852), .B1(n1637), .B2(n2863), .ZN(n2630)
         );
  OAI22_X1 U559 ( .A1(n1639), .A2(n2896), .B1(n1640), .B2(n2907), .ZN(n2631)
         );
  OAI22_X1 U560 ( .A1(n1599), .A2(n2852), .B1(n1600), .B2(n2863), .ZN(n2605)
         );
  OAI22_X1 U561 ( .A1(n1602), .A2(n2896), .B1(n1603), .B2(n2907), .ZN(n2606)
         );
  OAI22_X1 U562 ( .A1(n1562), .A2(n2851), .B1(n1563), .B2(n2862), .ZN(n2580)
         );
  OAI22_X1 U563 ( .A1(n1565), .A2(n2895), .B1(n1566), .B2(n2906), .ZN(n2581)
         );
  OAI22_X1 U564 ( .A1(n1525), .A2(n2852), .B1(n1526), .B2(n2863), .ZN(n2555)
         );
  OAI22_X1 U565 ( .A1(n1528), .A2(n2896), .B1(n1529), .B2(n2907), .ZN(n2556)
         );
  OAI22_X1 U566 ( .A1(n1488), .A2(n2853), .B1(n1489), .B2(n2864), .ZN(n2530)
         );
  OAI22_X1 U567 ( .A1(n1491), .A2(n2897), .B1(n1492), .B2(n2908), .ZN(n2531)
         );
  OAI22_X1 U568 ( .A1(n1414), .A2(n2853), .B1(n1415), .B2(n2864), .ZN(n2480)
         );
  OAI22_X1 U569 ( .A1(n1417), .A2(n2897), .B1(n1418), .B2(n2908), .ZN(n2481)
         );
  OAI22_X1 U570 ( .A1(n1377), .A2(n2852), .B1(n1378), .B2(n2863), .ZN(n2455)
         );
  OAI22_X1 U571 ( .A1(n1380), .A2(n2896), .B1(n1381), .B2(n2907), .ZN(n2456)
         );
  OAI22_X1 U572 ( .A1(n1340), .A2(n2852), .B1(n1341), .B2(n2863), .ZN(n2430)
         );
  OAI22_X1 U573 ( .A1(n1343), .A2(n2896), .B1(n1344), .B2(n2908), .ZN(n2431)
         );
  OAI22_X1 U574 ( .A1(n1303), .A2(n2852), .B1(n1304), .B2(n2863), .ZN(n2405)
         );
  OAI22_X1 U575 ( .A1(n1306), .A2(n2896), .B1(n1307), .B2(n2907), .ZN(n2406)
         );
  OAI22_X1 U576 ( .A1(n1266), .A2(n2853), .B1(n1267), .B2(n2864), .ZN(n2380)
         );
  OAI22_X1 U577 ( .A1(n1269), .A2(n2897), .B1(n1270), .B2(n2908), .ZN(n2381)
         );
  OAI22_X1 U578 ( .A1(n1229), .A2(n2853), .B1(n1230), .B2(n2864), .ZN(n2350)
         );
  OAI22_X1 U579 ( .A1(n1232), .A2(n2897), .B1(n1233), .B2(n2907), .ZN(n2351)
         );
  OAI22_X1 U580 ( .A1(n1192), .A2(n2853), .B1(n1193), .B2(n2864), .ZN(n2316)
         );
  OAI22_X1 U581 ( .A1(n1195), .A2(n2897), .B1(n1196), .B2(n2908), .ZN(n2318)
         );
  OAI22_X1 U582 ( .A1(n1155), .A2(n2852), .B1(n1156), .B2(n2863), .ZN(n2283)
         );
  OAI22_X1 U583 ( .A1(n1158), .A2(n2896), .B1(n1159), .B2(n2906), .ZN(n2284)
         );
  OAI22_X1 U584 ( .A1(n1118), .A2(n2853), .B1(n1119), .B2(n2864), .ZN(n2250)
         );
  OAI22_X1 U585 ( .A1(n1121), .A2(n2897), .B1(n1122), .B2(n2908), .ZN(n2251)
         );
  OAI22_X1 U586 ( .A1(n1081), .A2(n2852), .B1(n1082), .B2(n2863), .ZN(n2213)
         );
  OAI22_X1 U587 ( .A1(n1084), .A2(n2896), .B1(n1085), .B2(n2907), .ZN(n2214)
         );
  OAI22_X1 U588 ( .A1(n1007), .A2(n2853), .B1(n1008), .B2(n2864), .ZN(n2142)
         );
  OAI22_X1 U589 ( .A1(n1010), .A2(n2897), .B1(n1011), .B2(n2908), .ZN(n2143)
         );
  OAI22_X1 U590 ( .A1(n970), .A2(n2852), .B1(n971), .B2(n2863), .ZN(n2117) );
  OAI22_X1 U591 ( .A1(n973), .A2(n2896), .B1(n974), .B2(n2907), .ZN(n2118) );
  OAI22_X1 U592 ( .A1(n2978), .A2(n1902), .B1(n2967), .B2(n1903), .ZN(n1889)
         );
  OAI22_X1 U593 ( .A1(n2977), .A2(n1876), .B1(n2966), .B2(n1877), .ZN(n1868)
         );
  OAI22_X1 U594 ( .A1(n2983), .A2(n1474), .B1(n2972), .B2(n1475), .ZN(n1466)
         );
  OAI22_X1 U595 ( .A1(n2983), .A2(n1464), .B1(n2972), .B2(n1465), .ZN(n1456)
         );
  OAI22_X1 U596 ( .A1(n2980), .A2(n1067), .B1(n2969), .B2(n1068), .ZN(n1059)
         );
  OAI22_X1 U597 ( .A1(n2980), .A2(n1057), .B1(n2969), .B2(n1058), .ZN(n1049)
         );
  OAI22_X1 U598 ( .A1(n2979), .A2(n956), .B1(n2968), .B2(n957), .ZN(n948) );
  OAI22_X1 U599 ( .A1(n2979), .A2(n946), .B1(n2968), .B2(n947), .ZN(n938) );
  OAI22_X1 U600 ( .A1(n2979), .A2(n919), .B1(n2968), .B2(n920), .ZN(n911) );
  OAI22_X1 U601 ( .A1(n2979), .A2(n909), .B1(n2968), .B2(n910), .ZN(n901) );
  OAI22_X1 U602 ( .A1(n2979), .A2(n882), .B1(n2968), .B2(n883), .ZN(n874) );
  OAI22_X1 U603 ( .A1(n2979), .A2(n872), .B1(n2968), .B2(n873), .ZN(n864) );
  OAI22_X1 U604 ( .A1(n2979), .A2(n845), .B1(n2968), .B2(n846), .ZN(n837) );
  OAI22_X1 U605 ( .A1(n2978), .A2(n835), .B1(n2967), .B2(n836), .ZN(n827) );
  OAI22_X1 U606 ( .A1(n2978), .A2(n798), .B1(n2967), .B2(n799), .ZN(n790) );
  OAI22_X1 U607 ( .A1(n2978), .A2(n808), .B1(n2967), .B2(n809), .ZN(n800) );
  OAI22_X1 U608 ( .A1(n2978), .A2(n771), .B1(n2967), .B2(n772), .ZN(n763) );
  OAI22_X1 U609 ( .A1(n2978), .A2(n761), .B1(n2967), .B2(n762), .ZN(n753) );
  OAI22_X1 U610 ( .A1(n2978), .A2(n734), .B1(n2967), .B2(n735), .ZN(n726) );
  OAI22_X1 U611 ( .A1(n2978), .A2(n724), .B1(n2967), .B2(n725), .ZN(n716) );
  OAI22_X1 U612 ( .A1(n2985), .A2(n1834), .B1(n2974), .B2(n1835), .ZN(n1826)
         );
  OAI22_X1 U613 ( .A1(n2985), .A2(n1844), .B1(n2974), .B2(n1845), .ZN(n1836)
         );
  OAI22_X1 U614 ( .A1(n2985), .A2(n1807), .B1(n2974), .B2(n1808), .ZN(n1799)
         );
  OAI22_X1 U615 ( .A1(n2985), .A2(n1797), .B1(n2974), .B2(n1798), .ZN(n1789)
         );
  OAI22_X1 U616 ( .A1(n2985), .A2(n1770), .B1(n2974), .B2(n1771), .ZN(n1762)
         );
  OAI22_X1 U617 ( .A1(n2985), .A2(n1760), .B1(n2974), .B2(n1761), .ZN(n1752)
         );
  OAI22_X1 U618 ( .A1(n2985), .A2(n1723), .B1(n2974), .B2(n1724), .ZN(n1715)
         );
  OAI22_X1 U619 ( .A1(n2985), .A2(n1733), .B1(n2974), .B2(n1734), .ZN(n1725)
         );
  OAI22_X1 U620 ( .A1(n2984), .A2(n1696), .B1(n2973), .B2(n1697), .ZN(n1688)
         );
  OAI22_X1 U621 ( .A1(n2984), .A2(n1686), .B1(n2973), .B2(n1687), .ZN(n1678)
         );
  OAI22_X1 U622 ( .A1(n2984), .A2(n1659), .B1(n2973), .B2(n1660), .ZN(n1651)
         );
  OAI22_X1 U623 ( .A1(n2984), .A2(n1649), .B1(n2973), .B2(n1650), .ZN(n1641)
         );
  OAI22_X1 U624 ( .A1(n2984), .A2(n1622), .B1(n2973), .B2(n1623), .ZN(n1614)
         );
  OAI22_X1 U625 ( .A1(n2984), .A2(n1612), .B1(n2973), .B2(n1613), .ZN(n1604)
         );
  OAI22_X1 U626 ( .A1(n2984), .A2(n1585), .B1(n2973), .B2(n1586), .ZN(n1577)
         );
  OAI22_X1 U627 ( .A1(n2984), .A2(n1575), .B1(n2973), .B2(n1576), .ZN(n1567)
         );
  OAI22_X1 U628 ( .A1(n2983), .A2(n1548), .B1(n2972), .B2(n1549), .ZN(n1540)
         );
  OAI22_X1 U629 ( .A1(n2983), .A2(n1538), .B1(n2972), .B2(n1539), .ZN(n1530)
         );
  OAI22_X1 U630 ( .A1(n2983), .A2(n1511), .B1(n2972), .B2(n1512), .ZN(n1503)
         );
  OAI22_X1 U631 ( .A1(n2983), .A2(n1501), .B1(n2972), .B2(n1502), .ZN(n1493)
         );
  OAI22_X1 U632 ( .A1(n2983), .A2(n1437), .B1(n2972), .B2(n1438), .ZN(n1429)
         );
  OAI22_X1 U633 ( .A1(n2983), .A2(n1427), .B1(n2972), .B2(n1428), .ZN(n1419)
         );
  OAI22_X1 U634 ( .A1(n2982), .A2(n1400), .B1(n2971), .B2(n1401), .ZN(n1392)
         );
  OAI22_X1 U635 ( .A1(n2982), .A2(n1390), .B1(n2971), .B2(n1391), .ZN(n1382)
         );
  OAI22_X1 U636 ( .A1(n2982), .A2(n1363), .B1(n2971), .B2(n1364), .ZN(n1355)
         );
  OAI22_X1 U637 ( .A1(n2982), .A2(n1353), .B1(n2971), .B2(n1354), .ZN(n1345)
         );
  OAI22_X1 U638 ( .A1(n2982), .A2(n1326), .B1(n2971), .B2(n1327), .ZN(n1318)
         );
  OAI22_X1 U639 ( .A1(n2982), .A2(n1316), .B1(n2971), .B2(n1317), .ZN(n1308)
         );
  OAI22_X1 U640 ( .A1(n2982), .A2(n1289), .B1(n2971), .B2(n1290), .ZN(n1281)
         );
  OAI22_X1 U641 ( .A1(n2981), .A2(n1279), .B1(n2970), .B2(n1280), .ZN(n1271)
         );
  OAI22_X1 U642 ( .A1(n2981), .A2(n1252), .B1(n2970), .B2(n1253), .ZN(n1244)
         );
  OAI22_X1 U643 ( .A1(n2981), .A2(n1242), .B1(n2970), .B2(n1243), .ZN(n1234)
         );
  OAI22_X1 U644 ( .A1(n2981), .A2(n1215), .B1(n2970), .B2(n1216), .ZN(n1207)
         );
  OAI22_X1 U645 ( .A1(n2981), .A2(n1205), .B1(n2970), .B2(n1206), .ZN(n1197)
         );
  OAI22_X1 U646 ( .A1(n2981), .A2(n1178), .B1(n2970), .B2(n1179), .ZN(n1170)
         );
  OAI22_X1 U647 ( .A1(n2981), .A2(n1168), .B1(n2970), .B2(n1169), .ZN(n1160)
         );
  OAI22_X1 U648 ( .A1(n2981), .A2(n1141), .B1(n2970), .B2(n1142), .ZN(n1133)
         );
  OAI22_X1 U649 ( .A1(n2980), .A2(n1131), .B1(n2969), .B2(n1132), .ZN(n1123)
         );
  OAI22_X1 U650 ( .A1(n2980), .A2(n1104), .B1(n2969), .B2(n1105), .ZN(n1096)
         );
  OAI22_X1 U651 ( .A1(n2980), .A2(n1094), .B1(n2969), .B2(n1095), .ZN(n1086)
         );
  OAI22_X1 U652 ( .A1(n2980), .A2(n1030), .B1(n2969), .B2(n1031), .ZN(n1022)
         );
  OAI22_X1 U653 ( .A1(n2980), .A2(n1020), .B1(n2969), .B2(n1021), .ZN(n1012)
         );
  OAI22_X1 U654 ( .A1(n2980), .A2(n993), .B1(n2969), .B2(n994), .ZN(n985) );
  OAI22_X1 U655 ( .A1(n2979), .A2(n983), .B1(n2968), .B2(n984), .ZN(n975) );
  NOR2_X1 U656 ( .A1(n1854), .A2(read_address_2[0]), .ZN(n695) );
  NOR2_X1 U657 ( .A1(n1856), .A2(read_address_2[0]), .ZN(n697) );
  NOR2_X1 U658 ( .A1(n1857), .A2(read_address_2[0]), .ZN(n696) );
  BUF_X1 U659 ( .A(n687), .Z(n3031) );
  BUF_X1 U660 ( .A(n1928), .Z(n2822) );
  BUF_X1 U661 ( .A(n687), .Z(n3032) );
  NOR2_X1 U662 ( .A1(n1888), .A2(n1895), .ZN(n1899) );
  OAI21_X1 U663 ( .B1(n2764), .B2(n2765), .A(n2914), .ZN(n2763) );
  OAI221_X1 U664 ( .B1(n1903), .B2(n2869), .C1(n1902), .C2(n2850), .A(n2769), 
        .ZN(n2764) );
  OAI221_X1 U665 ( .B1(n1894), .B2(n2913), .C1(n1893), .C2(n2894), .A(n2768), 
        .ZN(n2765) );
  NOR2_X1 U666 ( .A1(n2785), .A2(n2786), .ZN(n2788) );
  NAND2_X1 U667 ( .A1(n2839), .A2(n3241), .ZN(n1941) );
  NAND2_X1 U668 ( .A1(n2875), .A2(n3241), .ZN(n1932) );
  NAND2_X1 U669 ( .A1(n2883), .A2(n3241), .ZN(n1930) );
  NAND2_X1 U670 ( .A1(n2831), .A2(n3241), .ZN(n1943) );
  AND2_X1 U671 ( .A1(n2766), .A2(n3240), .ZN(n1923) );
  AND2_X1 U672 ( .A1(n2766), .A2(n3241), .ZN(n1910) );
  NAND2_X1 U673 ( .A1(n1899), .A2(n1896), .ZN(n1855) );
  NAND2_X1 U674 ( .A1(n1901), .A2(n1896), .ZN(n707) );
  NAND2_X1 U675 ( .A1(n1898), .A2(n1896), .ZN(n705) );
  NAND2_X1 U676 ( .A1(n2789), .A2(n2787), .ZN(n1917) );
  NAND2_X1 U677 ( .A1(n2793), .A2(n2787), .ZN(n1916) );
  INV_X1 U678 ( .A(n1856), .ZN(n710) );
  INV_X1 U679 ( .A(n1857), .ZN(n709) );
  INV_X1 U680 ( .A(n1854), .ZN(n703) );
  AND2_X1 U681 ( .A1(n2788), .A2(n2787), .ZN(n1919) );
  OAI21_X1 U682 ( .B1(n662), .B2(n663), .A(n3044), .ZN(n2369) );
  OAI21_X1 U683 ( .B1(n662), .B2(n665), .A(n3044), .ZN(n2365) );
  OAI21_X1 U684 ( .B1(n662), .B2(n666), .A(n3044), .ZN(n2361) );
  OAI21_X1 U685 ( .B1(n662), .B2(n667), .A(n3044), .ZN(n2357) );
  OAI21_X1 U686 ( .B1(n662), .B2(n668), .A(n3044), .ZN(n2353) );
  OAI21_X1 U687 ( .B1(n662), .B2(n669), .A(n3044), .ZN(n2349) );
  OAI21_X1 U688 ( .B1(n662), .B2(n670), .A(n3044), .ZN(n2345) );
  OAI21_X1 U689 ( .B1(n662), .B2(n671), .A(n3044), .ZN(n2341) );
  OAI21_X1 U690 ( .B1(n663), .B2(n672), .A(n3044), .ZN(n2337) );
  OAI21_X1 U691 ( .B1(n665), .B2(n672), .A(n3044), .ZN(n2333) );
  OAI21_X1 U692 ( .B1(n666), .B2(n672), .A(n3044), .ZN(n2329) );
  OAI21_X1 U693 ( .B1(n667), .B2(n672), .A(n3044), .ZN(n2325) );
  OAI21_X1 U694 ( .B1(n668), .B2(n672), .A(n3045), .ZN(n2321) );
  OAI21_X1 U695 ( .B1(n669), .B2(n672), .A(n3045), .ZN(n2317) );
  OAI21_X1 U696 ( .B1(n670), .B2(n672), .A(n3045), .ZN(n2313) );
  OAI21_X1 U697 ( .B1(n671), .B2(n672), .A(n3045), .ZN(n2309) );
  OAI21_X1 U698 ( .B1(n663), .B2(n674), .A(n3045), .ZN(n2305) );
  OAI21_X1 U699 ( .B1(n665), .B2(n674), .A(n3045), .ZN(n2301) );
  OAI21_X1 U700 ( .B1(n666), .B2(n674), .A(n3045), .ZN(n2297) );
  OAI21_X1 U701 ( .B1(n667), .B2(n674), .A(n3045), .ZN(n2293) );
  OAI21_X1 U702 ( .B1(n668), .B2(n674), .A(n3045), .ZN(n2289) );
  OAI21_X1 U703 ( .B1(n669), .B2(n674), .A(n3045), .ZN(n2285) );
  OAI21_X1 U704 ( .B1(n670), .B2(n674), .A(n3045), .ZN(n2281) );
  OAI21_X1 U705 ( .B1(n671), .B2(n674), .A(n3045), .ZN(n2277) );
  OAI21_X1 U706 ( .B1(n663), .B2(n679), .A(n3046), .ZN(n2273) );
  OAI21_X1 U707 ( .B1(n665), .B2(n679), .A(n3046), .ZN(n2269) );
  OAI21_X1 U708 ( .B1(n666), .B2(n679), .A(n3046), .ZN(n2265) );
  OAI21_X1 U709 ( .B1(n667), .B2(n679), .A(n3046), .ZN(n2261) );
  OAI21_X1 U710 ( .B1(n668), .B2(n679), .A(n3046), .ZN(n2257) );
  OAI21_X1 U711 ( .B1(n669), .B2(n679), .A(n3046), .ZN(n2253) );
  OAI21_X1 U712 ( .B1(n670), .B2(n679), .A(n3046), .ZN(n2249) );
  BUF_X1 U713 ( .A(n2227), .Z(n3161) );
  BUF_X1 U714 ( .A(n2224), .Z(n3164) );
  BUF_X1 U715 ( .A(n2221), .Z(n3167) );
  BUF_X1 U716 ( .A(n2218), .Z(n3170) );
  BUF_X1 U717 ( .A(n2215), .Z(n3173) );
  BUF_X1 U718 ( .A(n2212), .Z(n3176) );
  BUF_X1 U719 ( .A(n2209), .Z(n3179) );
  BUF_X1 U720 ( .A(n2206), .Z(n3182) );
  BUF_X1 U721 ( .A(n2203), .Z(n3185) );
  BUF_X1 U722 ( .A(n2200), .Z(n3188) );
  BUF_X1 U723 ( .A(n2197), .Z(n3191) );
  BUF_X1 U724 ( .A(n2194), .Z(n3194) );
  BUF_X1 U725 ( .A(n2191), .Z(n3197) );
  BUF_X1 U726 ( .A(n2188), .Z(n3200) );
  BUF_X1 U727 ( .A(n2185), .Z(n3203) );
  BUF_X1 U728 ( .A(n2182), .Z(n3206) );
  BUF_X1 U729 ( .A(n2179), .Z(n3209) );
  BUF_X1 U730 ( .A(n2176), .Z(n3212) );
  BUF_X1 U731 ( .A(n2173), .Z(n3215) );
  BUF_X1 U732 ( .A(n2170), .Z(n3218) );
  BUF_X1 U733 ( .A(n2167), .Z(n3221) );
  BUF_X1 U734 ( .A(n2164), .Z(n3224) );
  BUF_X1 U735 ( .A(n2161), .Z(n3227) );
  BUF_X1 U736 ( .A(n2158), .Z(n3230) );
  BUF_X1 U737 ( .A(n2155), .Z(n3233) );
  BUF_X1 U738 ( .A(n2152), .Z(n3236) );
  BUF_X1 U739 ( .A(n2227), .Z(n3160) );
  BUF_X1 U740 ( .A(n2224), .Z(n3163) );
  BUF_X1 U741 ( .A(n2221), .Z(n3166) );
  BUF_X1 U742 ( .A(n2218), .Z(n3169) );
  BUF_X1 U743 ( .A(n2215), .Z(n3172) );
  BUF_X1 U744 ( .A(n2212), .Z(n3175) );
  BUF_X1 U745 ( .A(n2209), .Z(n3178) );
  BUF_X1 U746 ( .A(n2206), .Z(n3181) );
  BUF_X1 U747 ( .A(n2203), .Z(n3184) );
  BUF_X1 U748 ( .A(n2200), .Z(n3187) );
  BUF_X1 U749 ( .A(n2197), .Z(n3190) );
  BUF_X1 U750 ( .A(n2194), .Z(n3193) );
  BUF_X1 U751 ( .A(n2191), .Z(n3196) );
  BUF_X1 U752 ( .A(n2188), .Z(n3199) );
  BUF_X1 U753 ( .A(n2185), .Z(n3202) );
  BUF_X1 U754 ( .A(n2182), .Z(n3205) );
  BUF_X1 U755 ( .A(n2179), .Z(n3208) );
  BUF_X1 U756 ( .A(n2176), .Z(n3211) );
  BUF_X1 U757 ( .A(n2173), .Z(n3214) );
  BUF_X1 U758 ( .A(n2170), .Z(n3217) );
  BUF_X1 U759 ( .A(n2167), .Z(n3220) );
  BUF_X1 U760 ( .A(n2164), .Z(n3223) );
  BUF_X1 U761 ( .A(n2161), .Z(n3226) );
  BUF_X1 U762 ( .A(n2158), .Z(n3229) );
  BUF_X1 U763 ( .A(n2155), .Z(n3232) );
  BUF_X1 U764 ( .A(n2152), .Z(n3235) );
  BUF_X1 U765 ( .A(n2245), .Z(n3143) );
  BUF_X1 U766 ( .A(n2242), .Z(n3146) );
  BUF_X1 U767 ( .A(n2239), .Z(n3149) );
  BUF_X1 U768 ( .A(n2236), .Z(n3152) );
  BUF_X1 U769 ( .A(n2233), .Z(n3155) );
  BUF_X1 U770 ( .A(n2230), .Z(n3158) );
  BUF_X1 U771 ( .A(n2245), .Z(n3142) );
  BUF_X1 U772 ( .A(n2242), .Z(n3145) );
  BUF_X1 U773 ( .A(n2239), .Z(n3148) );
  BUF_X1 U774 ( .A(n2236), .Z(n3151) );
  BUF_X1 U775 ( .A(n2233), .Z(n3154) );
  BUF_X1 U776 ( .A(n2230), .Z(n3157) );
  BUF_X1 U777 ( .A(n2227), .Z(n3162) );
  BUF_X1 U778 ( .A(n2224), .Z(n3165) );
  BUF_X1 U779 ( .A(n2221), .Z(n3168) );
  BUF_X1 U780 ( .A(n2218), .Z(n3171) );
  BUF_X1 U781 ( .A(n2215), .Z(n3174) );
  BUF_X1 U782 ( .A(n2212), .Z(n3177) );
  BUF_X1 U783 ( .A(n2209), .Z(n3180) );
  BUF_X1 U784 ( .A(n2206), .Z(n3183) );
  BUF_X1 U785 ( .A(n2203), .Z(n3186) );
  BUF_X1 U786 ( .A(n2200), .Z(n3189) );
  BUF_X1 U787 ( .A(n2197), .Z(n3192) );
  BUF_X1 U788 ( .A(n2194), .Z(n3195) );
  BUF_X1 U789 ( .A(n2191), .Z(n3198) );
  BUF_X1 U790 ( .A(n2188), .Z(n3201) );
  BUF_X1 U791 ( .A(n2185), .Z(n3204) );
  BUF_X1 U792 ( .A(n2182), .Z(n3207) );
  BUF_X1 U793 ( .A(n2179), .Z(n3210) );
  BUF_X1 U794 ( .A(n2176), .Z(n3213) );
  BUF_X1 U795 ( .A(n2173), .Z(n3216) );
  BUF_X1 U796 ( .A(n2170), .Z(n3219) );
  BUF_X1 U797 ( .A(n2167), .Z(n3222) );
  BUF_X1 U798 ( .A(n2164), .Z(n3225) );
  BUF_X1 U799 ( .A(n2161), .Z(n3228) );
  BUF_X1 U800 ( .A(n2158), .Z(n3231) );
  BUF_X1 U801 ( .A(n2155), .Z(n3234) );
  BUF_X1 U802 ( .A(n2152), .Z(n3237) );
  BUF_X1 U803 ( .A(n2245), .Z(n3144) );
  BUF_X1 U804 ( .A(n2242), .Z(n3147) );
  BUF_X1 U805 ( .A(n2239), .Z(n3150) );
  BUF_X1 U806 ( .A(n2236), .Z(n3153) );
  BUF_X1 U807 ( .A(n2233), .Z(n3156) );
  BUF_X1 U808 ( .A(n2230), .Z(n3159) );
  BUF_X1 U809 ( .A(n664), .Z(n3042) );
  BUF_X1 U810 ( .A(n664), .Z(n3043) );
  NOR4_X1 U811 ( .A1(n2917), .A2(n1885), .A3(n1886), .A4(n1887), .ZN(n1883) );
  AOI22_X1 U812 ( .A1(n3035), .A2(n924), .B1(n3032), .B2(write_data[3]), .ZN(
        n923) );
  NAND4_X1 U813 ( .A1(n925), .A2(n926), .A3(n927), .A4(n928), .ZN(n924) );
  AOI22_X1 U814 ( .A1(\bank_register[20][3] ), .A2(n3017), .B1(
        \bank_register[28][3] ), .B2(n3014), .ZN(n926) );
  AOI22_X1 U815 ( .A1(\bank_register[24][3] ), .A2(n3023), .B1(
        \bank_register[12][3] ), .B2(n3020), .ZN(n927) );
  AOI22_X1 U816 ( .A1(n3035), .A2(n887), .B1(n3032), .B2(write_data[4]), .ZN(
        n886) );
  NAND4_X1 U817 ( .A1(n888), .A2(n889), .A3(n890), .A4(n891), .ZN(n887) );
  AOI22_X1 U818 ( .A1(\bank_register[20][4] ), .A2(n3017), .B1(
        \bank_register[28][4] ), .B2(n3014), .ZN(n889) );
  AOI22_X1 U819 ( .A1(\bank_register[24][4] ), .A2(n3023), .B1(
        \bank_register[12][4] ), .B2(n3020), .ZN(n890) );
  AOI22_X1 U820 ( .A1(n3035), .A2(n850), .B1(n3032), .B2(write_data[5]), .ZN(
        n849) );
  NAND4_X1 U821 ( .A1(n851), .A2(n852), .A3(n853), .A4(n854), .ZN(n850) );
  AOI22_X1 U822 ( .A1(\bank_register[20][5] ), .A2(n3017), .B1(
        \bank_register[28][5] ), .B2(n3014), .ZN(n852) );
  AOI22_X1 U823 ( .A1(\bank_register[24][5] ), .A2(n3023), .B1(
        \bank_register[12][5] ), .B2(n3020), .ZN(n853) );
  AOI22_X1 U824 ( .A1(n3035), .A2(n813), .B1(n3032), .B2(write_data[6]), .ZN(
        n812) );
  NAND4_X1 U825 ( .A1(n814), .A2(n815), .A3(n816), .A4(n817), .ZN(n813) );
  AOI22_X1 U826 ( .A1(\bank_register[20][6] ), .A2(n3017), .B1(
        \bank_register[28][6] ), .B2(n3014), .ZN(n815) );
  AOI22_X1 U827 ( .A1(\bank_register[24][6] ), .A2(n3023), .B1(
        \bank_register[12][6] ), .B2(n3020), .ZN(n816) );
  AOI22_X1 U828 ( .A1(n3035), .A2(n776), .B1(n3032), .B2(write_data[7]), .ZN(
        n775) );
  NAND4_X1 U829 ( .A1(n777), .A2(n778), .A3(n779), .A4(n780), .ZN(n776) );
  AOI22_X1 U830 ( .A1(\bank_register[20][7] ), .A2(n3017), .B1(
        \bank_register[28][7] ), .B2(n3014), .ZN(n778) );
  AOI22_X1 U831 ( .A1(\bank_register[24][7] ), .A2(n3023), .B1(
        \bank_register[12][7] ), .B2(n3020), .ZN(n779) );
  AOI22_X1 U832 ( .A1(n3035), .A2(n739), .B1(n3032), .B2(write_data[8]), .ZN(
        n738) );
  NAND4_X1 U833 ( .A1(n740), .A2(n741), .A3(n742), .A4(n743), .ZN(n739) );
  AOI22_X1 U834 ( .A1(\bank_register[20][8] ), .A2(n3017), .B1(
        \bank_register[28][8] ), .B2(n3014), .ZN(n741) );
  AOI22_X1 U835 ( .A1(\bank_register[24][8] ), .A2(n3023), .B1(
        \bank_register[12][8] ), .B2(n3020), .ZN(n742) );
  AOI22_X1 U836 ( .A1(n3035), .A2(n686), .B1(n3032), .B2(write_data[9]), .ZN(
        n684) );
  NAND4_X1 U837 ( .A1(n688), .A2(n689), .A3(n690), .A4(n691), .ZN(n686) );
  AOI22_X1 U838 ( .A1(\bank_register[20][9] ), .A2(n3017), .B1(
        \bank_register[28][9] ), .B2(n3014), .ZN(n689) );
  AOI22_X1 U839 ( .A1(\bank_register[24][9] ), .A2(n3023), .B1(
        \bank_register[12][9] ), .B2(n3020), .ZN(n690) );
  AOI22_X1 U840 ( .A1(n3035), .A2(n961), .B1(n3032), .B2(write_data[31]), .ZN(
        n960) );
  NAND4_X1 U841 ( .A1(n962), .A2(n963), .A3(n964), .A4(n965), .ZN(n961) );
  AOI22_X1 U842 ( .A1(\bank_register[20][31] ), .A2(n3017), .B1(
        \bank_register[28][31] ), .B2(n3014), .ZN(n963) );
  AOI22_X1 U843 ( .A1(\bank_register[24][31] ), .A2(n3023), .B1(
        \bank_register[12][31] ), .B2(n3020), .ZN(n964) );
  AOI22_X1 U844 ( .A1(n3033), .A2(n1849), .B1(n3030), .B2(write_data[0]), .ZN(
        n1848) );
  NAND4_X1 U845 ( .A1(n1850), .A2(n1851), .A3(n1852), .A4(n1853), .ZN(n1849)
         );
  AOI22_X1 U846 ( .A1(\bank_register[20][0] ), .A2(n3015), .B1(
        \bank_register[28][0] ), .B2(n3012), .ZN(n1851) );
  AOI22_X1 U847 ( .A1(\bank_register[24][0] ), .A2(n3021), .B1(
        \bank_register[12][0] ), .B2(n3018), .ZN(n1852) );
  AOI22_X1 U848 ( .A1(n3033), .A2(n1442), .B1(n3031), .B2(write_data[1]), .ZN(
        n1441) );
  NAND4_X1 U849 ( .A1(n1443), .A2(n1444), .A3(n1445), .A4(n1446), .ZN(n1442)
         );
  AOI22_X1 U850 ( .A1(\bank_register[20][1] ), .A2(n3015), .B1(
        \bank_register[28][1] ), .B2(n3012), .ZN(n1444) );
  AOI22_X1 U851 ( .A1(\bank_register[24][1] ), .A2(n3021), .B1(
        \bank_register[12][1] ), .B2(n3018), .ZN(n1445) );
  AOI22_X1 U852 ( .A1(n3034), .A2(n1035), .B1(n3031), .B2(write_data[2]), .ZN(
        n1034) );
  NAND4_X1 U853 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035)
         );
  AOI22_X1 U854 ( .A1(\bank_register[20][2] ), .A2(n3016), .B1(
        \bank_register[28][2] ), .B2(n3013), .ZN(n1037) );
  AOI22_X1 U855 ( .A1(\bank_register[24][2] ), .A2(n3022), .B1(
        \bank_register[12][2] ), .B2(n3019), .ZN(n1038) );
  AOI22_X1 U856 ( .A1(n3033), .A2(n1812), .B1(n3030), .B2(write_data[10]), 
        .ZN(n1811) );
  NAND4_X1 U857 ( .A1(n1813), .A2(n1814), .A3(n1815), .A4(n1816), .ZN(n1812)
         );
  AOI22_X1 U858 ( .A1(\bank_register[20][10] ), .A2(n3015), .B1(
        \bank_register[28][10] ), .B2(n3012), .ZN(n1814) );
  AOI22_X1 U859 ( .A1(\bank_register[24][10] ), .A2(n3021), .B1(
        \bank_register[12][10] ), .B2(n3018), .ZN(n1815) );
  AOI22_X1 U860 ( .A1(n3033), .A2(n1775), .B1(n3030), .B2(write_data[11]), 
        .ZN(n1774) );
  NAND4_X1 U861 ( .A1(n1776), .A2(n1777), .A3(n1778), .A4(n1779), .ZN(n1775)
         );
  AOI22_X1 U862 ( .A1(\bank_register[20][11] ), .A2(n3015), .B1(
        \bank_register[28][11] ), .B2(n3012), .ZN(n1777) );
  AOI22_X1 U863 ( .A1(\bank_register[24][11] ), .A2(n3021), .B1(
        \bank_register[12][11] ), .B2(n3018), .ZN(n1778) );
  AOI22_X1 U864 ( .A1(n3033), .A2(n1738), .B1(n3030), .B2(write_data[12]), 
        .ZN(n1737) );
  NAND4_X1 U865 ( .A1(n1739), .A2(n1740), .A3(n1741), .A4(n1742), .ZN(n1738)
         );
  AOI22_X1 U866 ( .A1(\bank_register[20][12] ), .A2(n3015), .B1(
        \bank_register[28][12] ), .B2(n3012), .ZN(n1740) );
  AOI22_X1 U867 ( .A1(\bank_register[24][12] ), .A2(n3021), .B1(
        \bank_register[12][12] ), .B2(n3018), .ZN(n1741) );
  AOI22_X1 U868 ( .A1(n3033), .A2(n1701), .B1(n3030), .B2(write_data[13]), 
        .ZN(n1700) );
  NAND4_X1 U869 ( .A1(n1702), .A2(n1703), .A3(n1704), .A4(n1705), .ZN(n1701)
         );
  AOI22_X1 U870 ( .A1(\bank_register[20][13] ), .A2(n3015), .B1(
        \bank_register[28][13] ), .B2(n3012), .ZN(n1703) );
  AOI22_X1 U871 ( .A1(\bank_register[24][13] ), .A2(n3021), .B1(
        \bank_register[12][13] ), .B2(n3018), .ZN(n1704) );
  AOI22_X1 U872 ( .A1(n3033), .A2(n1664), .B1(n3030), .B2(write_data[14]), 
        .ZN(n1663) );
  NAND4_X1 U873 ( .A1(n1665), .A2(n1666), .A3(n1667), .A4(n1668), .ZN(n1664)
         );
  AOI22_X1 U874 ( .A1(\bank_register[20][14] ), .A2(n3015), .B1(
        \bank_register[28][14] ), .B2(n3012), .ZN(n1666) );
  AOI22_X1 U875 ( .A1(\bank_register[24][14] ), .A2(n3021), .B1(
        \bank_register[12][14] ), .B2(n3018), .ZN(n1667) );
  AOI22_X1 U876 ( .A1(n3033), .A2(n1627), .B1(n3030), .B2(write_data[15]), 
        .ZN(n1626) );
  NAND4_X1 U877 ( .A1(n1628), .A2(n1629), .A3(n1630), .A4(n1631), .ZN(n1627)
         );
  AOI22_X1 U878 ( .A1(\bank_register[20][15] ), .A2(n3015), .B1(
        \bank_register[28][15] ), .B2(n3012), .ZN(n1629) );
  AOI22_X1 U879 ( .A1(\bank_register[24][15] ), .A2(n3021), .B1(
        \bank_register[12][15] ), .B2(n3018), .ZN(n1630) );
  AOI22_X1 U880 ( .A1(n3033), .A2(n1590), .B1(n3030), .B2(write_data[16]), 
        .ZN(n1589) );
  NAND4_X1 U881 ( .A1(n1591), .A2(n1592), .A3(n1593), .A4(n1594), .ZN(n1590)
         );
  AOI22_X1 U882 ( .A1(\bank_register[20][16] ), .A2(n3015), .B1(
        \bank_register[28][16] ), .B2(n3012), .ZN(n1592) );
  AOI22_X1 U883 ( .A1(\bank_register[24][16] ), .A2(n3021), .B1(
        \bank_register[12][16] ), .B2(n3018), .ZN(n1593) );
  AOI22_X1 U884 ( .A1(n3033), .A2(n1553), .B1(n3030), .B2(write_data[17]), 
        .ZN(n1552) );
  NAND4_X1 U885 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .ZN(n1553)
         );
  AOI22_X1 U886 ( .A1(\bank_register[20][17] ), .A2(n3015), .B1(
        \bank_register[28][17] ), .B2(n3012), .ZN(n1555) );
  AOI22_X1 U887 ( .A1(\bank_register[24][17] ), .A2(n3021), .B1(
        \bank_register[12][17] ), .B2(n3018), .ZN(n1556) );
  AOI22_X1 U888 ( .A1(n3033), .A2(n1516), .B1(n3030), .B2(write_data[18]), 
        .ZN(n1515) );
  NAND4_X1 U889 ( .A1(n1517), .A2(n1518), .A3(n1519), .A4(n1520), .ZN(n1516)
         );
  AOI22_X1 U890 ( .A1(\bank_register[20][18] ), .A2(n3015), .B1(
        \bank_register[28][18] ), .B2(n3012), .ZN(n1518) );
  AOI22_X1 U891 ( .A1(\bank_register[24][18] ), .A2(n3021), .B1(
        \bank_register[12][18] ), .B2(n3018), .ZN(n1519) );
  AOI22_X1 U892 ( .A1(n3033), .A2(n1479), .B1(n3030), .B2(write_data[19]), 
        .ZN(n1478) );
  NAND4_X1 U893 ( .A1(n1480), .A2(n1481), .A3(n1482), .A4(n1483), .ZN(n1479)
         );
  AOI22_X1 U894 ( .A1(\bank_register[20][19] ), .A2(n3015), .B1(
        \bank_register[28][19] ), .B2(n3012), .ZN(n1481) );
  AOI22_X1 U895 ( .A1(\bank_register[24][19] ), .A2(n3021), .B1(
        \bank_register[12][19] ), .B2(n3018), .ZN(n1482) );
  AOI22_X1 U896 ( .A1(n3034), .A2(n1405), .B1(n3031), .B2(write_data[20]), 
        .ZN(n1404) );
  NAND4_X1 U897 ( .A1(n1406), .A2(n1407), .A3(n1408), .A4(n1409), .ZN(n1405)
         );
  AOI22_X1 U898 ( .A1(\bank_register[20][20] ), .A2(n3016), .B1(
        \bank_register[28][20] ), .B2(n3013), .ZN(n1407) );
  AOI22_X1 U899 ( .A1(\bank_register[24][20] ), .A2(n3022), .B1(
        \bank_register[12][20] ), .B2(n3019), .ZN(n1408) );
  AOI22_X1 U900 ( .A1(n3034), .A2(n1368), .B1(n3031), .B2(write_data[21]), 
        .ZN(n1367) );
  NAND4_X1 U901 ( .A1(n1369), .A2(n1370), .A3(n1371), .A4(n1372), .ZN(n1368)
         );
  AOI22_X1 U902 ( .A1(\bank_register[20][21] ), .A2(n3016), .B1(
        \bank_register[28][21] ), .B2(n3013), .ZN(n1370) );
  AOI22_X1 U903 ( .A1(\bank_register[24][21] ), .A2(n3022), .B1(
        \bank_register[12][21] ), .B2(n3019), .ZN(n1371) );
  AOI22_X1 U904 ( .A1(n3034), .A2(n1331), .B1(n3031), .B2(write_data[22]), 
        .ZN(n1330) );
  NAND4_X1 U905 ( .A1(n1332), .A2(n1333), .A3(n1334), .A4(n1335), .ZN(n1331)
         );
  AOI22_X1 U906 ( .A1(\bank_register[20][22] ), .A2(n3016), .B1(
        \bank_register[28][22] ), .B2(n3013), .ZN(n1333) );
  AOI22_X1 U907 ( .A1(\bank_register[24][22] ), .A2(n3022), .B1(
        \bank_register[12][22] ), .B2(n3019), .ZN(n1334) );
  AOI22_X1 U908 ( .A1(n3034), .A2(n1294), .B1(n3031), .B2(write_data[23]), 
        .ZN(n1293) );
  NAND4_X1 U909 ( .A1(n1295), .A2(n1296), .A3(n1297), .A4(n1298), .ZN(n1294)
         );
  AOI22_X1 U910 ( .A1(\bank_register[20][23] ), .A2(n3016), .B1(
        \bank_register[28][23] ), .B2(n3013), .ZN(n1296) );
  AOI22_X1 U911 ( .A1(\bank_register[24][23] ), .A2(n3022), .B1(
        \bank_register[12][23] ), .B2(n3019), .ZN(n1297) );
  AOI22_X1 U912 ( .A1(n3034), .A2(n1257), .B1(n3031), .B2(write_data[24]), 
        .ZN(n1256) );
  NAND4_X1 U913 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1257)
         );
  AOI22_X1 U914 ( .A1(\bank_register[20][24] ), .A2(n3016), .B1(
        \bank_register[28][24] ), .B2(n3013), .ZN(n1259) );
  AOI22_X1 U915 ( .A1(\bank_register[24][24] ), .A2(n3022), .B1(
        \bank_register[12][24] ), .B2(n3019), .ZN(n1260) );
  AOI22_X1 U916 ( .A1(n3034), .A2(n1220), .B1(n3031), .B2(write_data[25]), 
        .ZN(n1219) );
  NAND4_X1 U917 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220)
         );
  AOI22_X1 U918 ( .A1(\bank_register[20][25] ), .A2(n3016), .B1(
        \bank_register[28][25] ), .B2(n3013), .ZN(n1222) );
  AOI22_X1 U919 ( .A1(\bank_register[24][25] ), .A2(n3022), .B1(
        \bank_register[12][25] ), .B2(n3019), .ZN(n1223) );
  AOI22_X1 U920 ( .A1(n3034), .A2(n1183), .B1(n3031), .B2(write_data[26]), 
        .ZN(n1182) );
  NAND4_X1 U921 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183)
         );
  AOI22_X1 U922 ( .A1(\bank_register[20][26] ), .A2(n3016), .B1(
        \bank_register[28][26] ), .B2(n3013), .ZN(n1185) );
  AOI22_X1 U923 ( .A1(\bank_register[24][26] ), .A2(n3022), .B1(
        \bank_register[12][26] ), .B2(n3019), .ZN(n1186) );
  AOI22_X1 U924 ( .A1(n3034), .A2(n1146), .B1(n3031), .B2(write_data[27]), 
        .ZN(n1145) );
  NAND4_X1 U925 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146)
         );
  AOI22_X1 U926 ( .A1(\bank_register[20][27] ), .A2(n3016), .B1(
        \bank_register[28][27] ), .B2(n3013), .ZN(n1148) );
  AOI22_X1 U927 ( .A1(\bank_register[24][27] ), .A2(n3022), .B1(
        \bank_register[12][27] ), .B2(n3019), .ZN(n1149) );
  AOI22_X1 U928 ( .A1(n3034), .A2(n1109), .B1(n3031), .B2(write_data[28]), 
        .ZN(n1108) );
  NAND4_X1 U929 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1109)
         );
  AOI22_X1 U930 ( .A1(\bank_register[20][28] ), .A2(n3016), .B1(
        \bank_register[28][28] ), .B2(n3013), .ZN(n1111) );
  AOI22_X1 U931 ( .A1(\bank_register[24][28] ), .A2(n3022), .B1(
        \bank_register[12][28] ), .B2(n3019), .ZN(n1112) );
  AOI22_X1 U932 ( .A1(n3034), .A2(n1072), .B1(n3031), .B2(write_data[29]), 
        .ZN(n1071) );
  NAND4_X1 U933 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072)
         );
  AOI22_X1 U934 ( .A1(\bank_register[20][29] ), .A2(n3016), .B1(
        \bank_register[28][29] ), .B2(n3013), .ZN(n1074) );
  AOI22_X1 U935 ( .A1(\bank_register[24][29] ), .A2(n3022), .B1(
        \bank_register[12][29] ), .B2(n3019), .ZN(n1075) );
  AOI22_X1 U936 ( .A1(n3034), .A2(n998), .B1(n3031), .B2(write_data[30]), .ZN(
        n997) );
  NAND4_X1 U937 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(n998) );
  AOI22_X1 U938 ( .A1(\bank_register[20][30] ), .A2(n3016), .B1(
        \bank_register[28][30] ), .B2(n3013), .ZN(n1000) );
  AOI22_X1 U939 ( .A1(\bank_register[24][30] ), .A2(n3022), .B1(
        \bank_register[12][30] ), .B2(n3019), .ZN(n1001) );
  INV_X1 U940 ( .A(read_address_1[0]), .ZN(n3241) );
  NAND4_X1 U941 ( .A1(n2794), .A2(n2795), .A3(n2796), .A4(n2797), .ZN(n2772)
         );
  NOR3_X1 U942 ( .A1(n2798), .A2(n1885), .A3(n2799), .ZN(n2797) );
  NOR2_X1 U943 ( .A1(n3030), .A2(read_address_2[1]), .ZN(n685) );
  INV_X1 U944 ( .A(read_address_1[3]), .ZN(n2785) );
  INV_X1 U945 ( .A(reg_write), .ZN(n1885) );
  AND4_X1 U946 ( .A1(n1880), .A2(n1881), .A3(n1882), .A4(n1883), .ZN(n687) );
  OAI21_X1 U947 ( .B1(n2084), .B2(n2085), .A(n2822), .ZN(n2073) );
  OAI221_X1 U948 ( .B1(n2094), .B2(n2810), .C1(n2095), .C2(n2807), .A(n2096), 
        .ZN(n2084) );
  OAI221_X1 U949 ( .B1(n2086), .B2(n2819), .C1(n2087), .C2(n2816), .A(n2088), 
        .ZN(n2085) );
  INV_X1 U950 ( .A(\bank_register[12][3] ), .ZN(n2095) );
  OAI21_X1 U951 ( .B1(n2059), .B2(n2060), .A(n2822), .ZN(n2048) );
  OAI221_X1 U952 ( .B1(n2069), .B2(n2810), .C1(n2070), .C2(n2807), .A(n2071), 
        .ZN(n2059) );
  OAI221_X1 U953 ( .B1(n2061), .B2(n2819), .C1(n2062), .C2(n2816), .A(n2063), 
        .ZN(n2060) );
  INV_X1 U954 ( .A(\bank_register[12][4] ), .ZN(n2070) );
  OAI21_X1 U955 ( .B1(n2034), .B2(n2035), .A(n2822), .ZN(n2023) );
  OAI221_X1 U956 ( .B1(n2044), .B2(n2810), .C1(n2045), .C2(n2807), .A(n2046), 
        .ZN(n2034) );
  OAI221_X1 U957 ( .B1(n2036), .B2(n2819), .C1(n2037), .C2(n2816), .A(n2038), 
        .ZN(n2035) );
  INV_X1 U958 ( .A(\bank_register[12][5] ), .ZN(n2045) );
  OAI21_X1 U959 ( .B1(n2009), .B2(n2010), .A(n2822), .ZN(n1998) );
  OAI221_X1 U960 ( .B1(n2019), .B2(n2810), .C1(n2020), .C2(n2807), .A(n2021), 
        .ZN(n2009) );
  OAI221_X1 U961 ( .B1(n2011), .B2(n2819), .C1(n2012), .C2(n2816), .A(n2013), 
        .ZN(n2010) );
  INV_X1 U962 ( .A(\bank_register[12][6] ), .ZN(n2020) );
  OAI21_X1 U963 ( .B1(n1984), .B2(n1985), .A(n2822), .ZN(n1973) );
  OAI221_X1 U964 ( .B1(n1994), .B2(n2810), .C1(n1995), .C2(n2807), .A(n1996), 
        .ZN(n1984) );
  OAI221_X1 U965 ( .B1(n1986), .B2(n2819), .C1(n1987), .C2(n2816), .A(n1988), 
        .ZN(n1985) );
  INV_X1 U966 ( .A(\bank_register[12][7] ), .ZN(n1995) );
  OAI21_X1 U967 ( .B1(n1959), .B2(n1960), .A(n2822), .ZN(n1948) );
  OAI221_X1 U968 ( .B1(n1969), .B2(n2810), .C1(n1970), .C2(n2807), .A(n1971), 
        .ZN(n1959) );
  OAI221_X1 U969 ( .B1(n1961), .B2(n2819), .C1(n1962), .C2(n2816), .A(n1963), 
        .ZN(n1960) );
  INV_X1 U970 ( .A(\bank_register[12][8] ), .ZN(n1970) );
  OAI21_X1 U971 ( .B1(n1926), .B2(n1927), .A(n2822), .ZN(n1905) );
  OAI221_X1 U972 ( .B1(n1940), .B2(n2810), .C1(n1942), .C2(n2807), .A(n1944), 
        .ZN(n1926) );
  OAI221_X1 U973 ( .B1(n1929), .B2(n2819), .C1(n1931), .C2(n2816), .A(n1933), 
        .ZN(n1927) );
  INV_X1 U974 ( .A(\bank_register[12][9] ), .ZN(n1942) );
  OAI221_X1 U975 ( .B1(n1873), .B2(n2909), .C1(n1872), .C2(n2898), .A(n2773), 
        .ZN(n2771) );
  AOI22_X1 U976 ( .A1(n2891), .A2(\bank_register[23][0] ), .B1(n2876), .B2(
        \bank_register[31][0] ), .ZN(n2773) );
  OAI221_X1 U977 ( .B1(n1054), .B2(n2910), .C1(n1053), .C2(n2899), .A(n2160), 
        .ZN(n2159) );
  AOI22_X1 U978 ( .A1(n2888), .A2(\bank_register[23][2] ), .B1(n2877), .B2(
        \bank_register[31][2] ), .ZN(n2160) );
  OAI221_X1 U979 ( .B1(n943), .B2(n2909), .C1(n942), .C2(n2898), .A(n2082), 
        .ZN(n2081) );
  AOI22_X1 U980 ( .A1(n2887), .A2(\bank_register[23][3] ), .B1(n2876), .B2(
        \bank_register[31][3] ), .ZN(n2082) );
  OAI221_X1 U981 ( .B1(n906), .B2(n2909), .C1(n905), .C2(n2898), .A(n2057), 
        .ZN(n2056) );
  AOI22_X1 U982 ( .A1(n2888), .A2(\bank_register[23][4] ), .B1(n2876), .B2(
        \bank_register[31][4] ), .ZN(n2057) );
  OAI221_X1 U983 ( .B1(n869), .B2(n2908), .C1(n868), .C2(n2898), .A(n2032), 
        .ZN(n2031) );
  AOI22_X1 U984 ( .A1(n2887), .A2(\bank_register[23][5] ), .B1(n2876), .B2(
        \bank_register[31][5] ), .ZN(n2032) );
  OAI221_X1 U985 ( .B1(n832), .B2(n2908), .C1(n831), .C2(n2897), .A(n2007), 
        .ZN(n2006) );
  AOI22_X1 U986 ( .A1(n2887), .A2(\bank_register[23][6] ), .B1(n2875), .B2(
        \bank_register[31][6] ), .ZN(n2007) );
  OAI221_X1 U987 ( .B1(n795), .B2(n2909), .C1(n794), .C2(n2898), .A(n1982), 
        .ZN(n1981) );
  AOI22_X1 U988 ( .A1(n2886), .A2(\bank_register[23][7] ), .B1(n2876), .B2(
        \bank_register[31][7] ), .ZN(n1982) );
  OAI221_X1 U989 ( .B1(n758), .B2(n2910), .C1(n757), .C2(n2898), .A(n1957), 
        .ZN(n1956) );
  AOI22_X1 U990 ( .A1(n2886), .A2(\bank_register[23][8] ), .B1(n2876), .B2(
        \bank_register[31][8] ), .ZN(n1957) );
  OAI221_X1 U991 ( .B1(n721), .B2(n2909), .C1(n720), .C2(n2899), .A(n1924), 
        .ZN(n1922) );
  AOI22_X1 U992 ( .A1(n2887), .A2(\bank_register[23][9] ), .B1(n2877), .B2(
        \bank_register[31][9] ), .ZN(n1924) );
  OAI221_X1 U993 ( .B1(n1387), .B2(n2911), .C1(n1386), .C2(n2900), .A(n2445), 
        .ZN(n2444) );
  AOI22_X1 U994 ( .A1(n2889), .A2(\bank_register[23][21] ), .B1(n2878), .B2(
        \bank_register[31][21] ), .ZN(n2445) );
  OAI221_X1 U995 ( .B1(n1350), .B2(n2911), .C1(n1349), .C2(n2900), .A(n2420), 
        .ZN(n2419) );
  AOI22_X1 U996 ( .A1(n2889), .A2(\bank_register[23][22] ), .B1(n2878), .B2(
        \bank_register[31][22] ), .ZN(n2420) );
  OAI221_X1 U997 ( .B1(n1313), .B2(n2911), .C1(n1312), .C2(n2900), .A(n2395), 
        .ZN(n2394) );
  AOI22_X1 U998 ( .A1(n2889), .A2(\bank_register[23][23] ), .B1(n2878), .B2(
        \bank_register[31][23] ), .ZN(n2395) );
  OAI221_X1 U999 ( .B1(n1276), .B2(n2911), .C1(n1275), .C2(n2900), .A(n2370), 
        .ZN(n2368) );
  AOI22_X1 U1000 ( .A1(n2889), .A2(\bank_register[23][24] ), .B1(n2878), .B2(
        \bank_register[31][24] ), .ZN(n2370) );
  OAI221_X1 U1001 ( .B1(n1239), .B2(n2911), .C1(n1238), .C2(n2900), .A(n2336), 
        .ZN(n2335) );
  AOI22_X1 U1002 ( .A1(n2889), .A2(\bank_register[23][25] ), .B1(n2878), .B2(
        \bank_register[31][25] ), .ZN(n2336) );
  OAI221_X1 U1003 ( .B1(n1202), .B2(n2910), .C1(n1201), .C2(n2900), .A(n2303), 
        .ZN(n2302) );
  AOI22_X1 U1004 ( .A1(n2888), .A2(\bank_register[23][26] ), .B1(n2878), .B2(
        \bank_register[31][26] ), .ZN(n2303) );
  OAI221_X1 U1005 ( .B1(n1165), .B2(n2910), .C1(n1164), .C2(n2899), .A(n2270), 
        .ZN(n2268) );
  AOI22_X1 U1006 ( .A1(n2888), .A2(\bank_register[23][27] ), .B1(n2877), .B2(
        \bank_register[31][27] ), .ZN(n2270) );
  OAI221_X1 U1007 ( .B1(n1128), .B2(n2910), .C1(n1127), .C2(n2899), .A(n2235), 
        .ZN(n2234) );
  AOI22_X1 U1008 ( .A1(n2888), .A2(\bank_register[23][28] ), .B1(n2877), .B2(
        \bank_register[31][28] ), .ZN(n2235) );
  OAI221_X1 U1009 ( .B1(n1091), .B2(n2910), .C1(n1090), .C2(n2899), .A(n2198), 
        .ZN(n2196) );
  AOI22_X1 U1010 ( .A1(n2888), .A2(\bank_register[23][29] ), .B1(n2877), .B2(
        \bank_register[31][29] ), .ZN(n2198) );
  OAI221_X1 U1011 ( .B1(n1017), .B2(n2909), .C1(n1016), .C2(n2898), .A(n2132), 
        .ZN(n2131) );
  AOI22_X1 U1012 ( .A1(n2888), .A2(\bank_register[23][30] ), .B1(n2876), .B2(
        \bank_register[31][30] ), .ZN(n2132) );
  OAI221_X1 U1013 ( .B1(n980), .B2(n2909), .C1(n979), .C2(n2898), .A(n2107), 
        .ZN(n2106) );
  AOI22_X1 U1014 ( .A1(n2887), .A2(\bank_register[23][31] ), .B1(n2876), .B2(
        \bank_register[31][31] ), .ZN(n2107) );
  OAI221_X1 U1015 ( .B1(n836), .B2(n2864), .C1(n835), .C2(n2853), .A(n2008), 
        .ZN(n2005) );
  AOI22_X1 U1016 ( .A1(n2843), .A2(\bank_register[27][6] ), .B1(n2831), .B2(
        \bank_register[15][6] ), .ZN(n2008) );
  OAI221_X1 U1017 ( .B1(n1428), .B2(n2867), .C1(n1427), .C2(n2857), .A(n2471), 
        .ZN(n2468) );
  AOI22_X1 U1018 ( .A1(n2845), .A2(\bank_register[27][20] ), .B1(n2835), .B2(
        \bank_register[15][20] ), .ZN(n2471) );
  AOI22_X1 U1019 ( .A1(\bank_register[8][3] ), .A2(n3029), .B1(
        \bank_register[16][3] ), .B2(n3026), .ZN(n928) );
  AOI22_X1 U1020 ( .A1(\bank_register[8][4] ), .A2(n3029), .B1(
        \bank_register[16][4] ), .B2(n3026), .ZN(n891) );
  AOI22_X1 U1021 ( .A1(\bank_register[8][5] ), .A2(n3029), .B1(
        \bank_register[16][5] ), .B2(n3026), .ZN(n854) );
  AOI22_X1 U1022 ( .A1(\bank_register[8][6] ), .A2(n3029), .B1(
        \bank_register[16][6] ), .B2(n3026), .ZN(n817) );
  AOI22_X1 U1023 ( .A1(\bank_register[8][7] ), .A2(n3029), .B1(
        \bank_register[16][7] ), .B2(n3026), .ZN(n780) );
  AOI22_X1 U1024 ( .A1(\bank_register[8][8] ), .A2(n3029), .B1(
        \bank_register[16][8] ), .B2(n3026), .ZN(n743) );
  AOI22_X1 U1025 ( .A1(\bank_register[8][9] ), .A2(n3029), .B1(
        \bank_register[16][9] ), .B2(n3026), .ZN(n691) );
  AOI22_X1 U1026 ( .A1(\bank_register[8][31] ), .A2(n3029), .B1(
        \bank_register[16][31] ), .B2(n3026), .ZN(n965) );
  AOI22_X1 U1027 ( .A1(\bank_register[8][0] ), .A2(n3027), .B1(
        \bank_register[16][0] ), .B2(n3024), .ZN(n1853) );
  AOI22_X1 U1028 ( .A1(\bank_register[8][1] ), .A2(n3027), .B1(
        \bank_register[16][1] ), .B2(n3024), .ZN(n1446) );
  AOI22_X1 U1029 ( .A1(\bank_register[8][2] ), .A2(n3028), .B1(
        \bank_register[16][2] ), .B2(n3025), .ZN(n1039) );
  AOI22_X1 U1030 ( .A1(\bank_register[8][10] ), .A2(n3027), .B1(
        \bank_register[16][10] ), .B2(n3024), .ZN(n1816) );
  AOI22_X1 U1031 ( .A1(\bank_register[8][11] ), .A2(n3027), .B1(
        \bank_register[16][11] ), .B2(n3024), .ZN(n1779) );
  AOI22_X1 U1032 ( .A1(\bank_register[8][12] ), .A2(n3027), .B1(
        \bank_register[16][12] ), .B2(n3024), .ZN(n1742) );
  AOI22_X1 U1033 ( .A1(\bank_register[8][13] ), .A2(n3027), .B1(
        \bank_register[16][13] ), .B2(n3024), .ZN(n1705) );
  AOI22_X1 U1034 ( .A1(\bank_register[8][14] ), .A2(n3027), .B1(
        \bank_register[16][14] ), .B2(n3024), .ZN(n1668) );
  AOI22_X1 U1035 ( .A1(\bank_register[8][15] ), .A2(n3027), .B1(
        \bank_register[16][15] ), .B2(n3024), .ZN(n1631) );
  AOI22_X1 U1036 ( .A1(\bank_register[8][16] ), .A2(n3027), .B1(
        \bank_register[16][16] ), .B2(n3024), .ZN(n1594) );
  AOI22_X1 U1037 ( .A1(\bank_register[8][17] ), .A2(n3027), .B1(
        \bank_register[16][17] ), .B2(n3024), .ZN(n1557) );
  AOI22_X1 U1038 ( .A1(\bank_register[8][18] ), .A2(n3027), .B1(
        \bank_register[16][18] ), .B2(n3024), .ZN(n1520) );
  AOI22_X1 U1039 ( .A1(\bank_register[8][19] ), .A2(n3027), .B1(
        \bank_register[16][19] ), .B2(n3024), .ZN(n1483) );
  AOI22_X1 U1040 ( .A1(\bank_register[8][20] ), .A2(n3028), .B1(
        \bank_register[16][20] ), .B2(n3025), .ZN(n1409) );
  AOI22_X1 U1041 ( .A1(\bank_register[8][21] ), .A2(n3028), .B1(
        \bank_register[16][21] ), .B2(n3025), .ZN(n1372) );
  AOI22_X1 U1042 ( .A1(\bank_register[8][22] ), .A2(n3028), .B1(
        \bank_register[16][22] ), .B2(n3025), .ZN(n1335) );
  AOI22_X1 U1043 ( .A1(\bank_register[8][23] ), .A2(n3028), .B1(
        \bank_register[16][23] ), .B2(n3025), .ZN(n1298) );
  AOI22_X1 U1044 ( .A1(\bank_register[8][24] ), .A2(n3028), .B1(
        \bank_register[16][24] ), .B2(n3025), .ZN(n1261) );
  AOI22_X1 U1045 ( .A1(\bank_register[8][25] ), .A2(n3028), .B1(
        \bank_register[16][25] ), .B2(n3025), .ZN(n1224) );
  AOI22_X1 U1046 ( .A1(\bank_register[8][26] ), .A2(n3028), .B1(
        \bank_register[16][26] ), .B2(n3025), .ZN(n1187) );
  AOI22_X1 U1047 ( .A1(\bank_register[8][27] ), .A2(n3028), .B1(
        \bank_register[16][27] ), .B2(n3025), .ZN(n1150) );
  AOI22_X1 U1048 ( .A1(\bank_register[8][28] ), .A2(n3028), .B1(
        \bank_register[16][28] ), .B2(n3025), .ZN(n1113) );
  AOI22_X1 U1049 ( .A1(\bank_register[8][29] ), .A2(n3028), .B1(
        \bank_register[16][29] ), .B2(n3025), .ZN(n1076) );
  AOI22_X1 U1050 ( .A1(\bank_register[8][30] ), .A2(n3028), .B1(
        \bank_register[16][30] ), .B2(n3025), .ZN(n1002) );
  AOI22_X1 U1051 ( .A1(n2811), .A2(\bank_register[4][0] ), .B1(
        read_address_1[0]), .B2(n2780), .ZN(n2779) );
  NAND2_X1 U1052 ( .A1(n2781), .A2(n2782), .ZN(n2780) );
  AOI221_X1 U1053 ( .B1(n2884), .B2(\bank_register[21][0] ), .C1(n2873), .C2(
        \bank_register[29][0] ), .A(n2784), .ZN(n2781) );
  AOI221_X1 U1054 ( .B1(n2840), .B2(\bank_register[25][0] ), .C1(n2829), .C2(
        \bank_register[13][0] ), .A(n2783), .ZN(n2782) );
  AOI22_X1 U1055 ( .A1(n2802), .A2(\bank_register[8][0] ), .B1(n2767), .B2(
        \bank_register[16][0] ), .ZN(n2792) );
  AOI22_X1 U1056 ( .A1(n2891), .A2(\bank_register[22][0] ), .B1(n2872), .B2(
        \bank_register[30][0] ), .ZN(n2768) );
  AOI22_X1 U1057 ( .A1(n2847), .A2(\bank_register[26][0] ), .B1(n2828), .B2(
        \bank_register[14][0] ), .ZN(n2769) );
  AOI22_X1 U1058 ( .A1(n2811), .A2(\bank_register[4][1] ), .B1(
        read_address_1[0]), .B2(n2502), .ZN(n2501) );
  NAND2_X1 U1059 ( .A1(n2503), .A2(n2504), .ZN(n2502) );
  AOI221_X1 U1060 ( .B1(n2884), .B2(\bank_register[21][1] ), .C1(n2874), .C2(
        \bank_register[29][1] ), .A(n2506), .ZN(n2503) );
  AOI221_X1 U1061 ( .B1(n2840), .B2(\bank_register[25][1] ), .C1(n2830), .C2(
        \bank_register[13][1] ), .A(n2505), .ZN(n2504) );
  AOI22_X1 U1062 ( .A1(n2802), .A2(\bank_register[8][1] ), .B1(n2767), .B2(
        \bank_register[16][1] ), .ZN(n2509) );
  AOI22_X1 U1063 ( .A1(n2890), .A2(\bank_register[22][1] ), .B1(n2879), .B2(
        \bank_register[30][1] ), .ZN(n2491) );
  AOI22_X1 U1064 ( .A1(n2812), .A2(\bank_register[4][2] ), .B1(
        read_address_1[0]), .B2(n2171), .ZN(n2169) );
  NAND2_X1 U1065 ( .A1(n2172), .A2(n2174), .ZN(n2171) );
  AOI221_X1 U1066 ( .B1(n2885), .B2(\bank_register[21][2] ), .C1(n2875), .C2(
        \bank_register[29][2] ), .A(n2177), .ZN(n2172) );
  AOI221_X1 U1067 ( .B1(n2841), .B2(\bank_register[25][2] ), .C1(n2831), .C2(
        \bank_register[13][2] ), .A(n2175), .ZN(n2174) );
  AOI22_X1 U1068 ( .A1(n2803), .A2(\bank_register[8][2] ), .B1(n2800), .B2(
        \bank_register[16][2] ), .ZN(n2181) );
  AOI22_X1 U1069 ( .A1(n2887), .A2(\bank_register[22][2] ), .B1(n2877), .B2(
        \bank_register[30][2] ), .ZN(n2154) );
  AOI22_X1 U1070 ( .A1(n2813), .A2(\bank_register[4][3] ), .B1(n3240), .B2(
        n2089), .ZN(n2088) );
  NAND2_X1 U1071 ( .A1(n2090), .A2(n2091), .ZN(n2089) );
  AOI221_X1 U1072 ( .B1(n2886), .B2(\bank_register[21][3] ), .C1(n2873), .C2(
        \bank_register[29][3] ), .A(n2093), .ZN(n2090) );
  AOI221_X1 U1073 ( .B1(n2842), .B2(\bank_register[25][3] ), .C1(n2829), .C2(
        \bank_register[13][3] ), .A(n2092), .ZN(n2091) );
  AOI22_X1 U1074 ( .A1(n2804), .A2(\bank_register[8][3] ), .B1(n2801), .B2(
        \bank_register[16][3] ), .ZN(n2096) );
  AOI22_X1 U1075 ( .A1(n2887), .A2(\bank_register[22][3] ), .B1(n2876), .B2(
        \bank_register[30][3] ), .ZN(n2078) );
  AOI22_X1 U1076 ( .A1(n2813), .A2(\bank_register[4][4] ), .B1(
        read_address_1[0]), .B2(n2064), .ZN(n2063) );
  NAND2_X1 U1077 ( .A1(n2065), .A2(n2066), .ZN(n2064) );
  AOI221_X1 U1078 ( .B1(n2885), .B2(\bank_register[21][4] ), .C1(n2874), .C2(
        \bank_register[29][4] ), .A(n2068), .ZN(n2065) );
  AOI221_X1 U1079 ( .B1(n2841), .B2(\bank_register[25][4] ), .C1(n2830), .C2(
        \bank_register[13][4] ), .A(n2067), .ZN(n2066) );
  AOI22_X1 U1080 ( .A1(n2804), .A2(\bank_register[8][4] ), .B1(n2801), .B2(
        \bank_register[16][4] ), .ZN(n2071) );
  AOI22_X1 U1081 ( .A1(n2887), .A2(\bank_register[22][4] ), .B1(n2876), .B2(
        \bank_register[30][4] ), .ZN(n2053) );
  AOI22_X1 U1082 ( .A1(n2813), .A2(\bank_register[4][5] ), .B1(
        read_address_1[0]), .B2(n2039), .ZN(n2038) );
  NAND2_X1 U1083 ( .A1(n2040), .A2(n2041), .ZN(n2039) );
  AOI221_X1 U1084 ( .B1(n2884), .B2(\bank_register[21][5] ), .C1(n2873), .C2(
        \bank_register[29][5] ), .A(n2043), .ZN(n2040) );
  AOI221_X1 U1085 ( .B1(n2840), .B2(\bank_register[25][5] ), .C1(n2829), .C2(
        \bank_register[13][5] ), .A(n2042), .ZN(n2041) );
  AOI22_X1 U1086 ( .A1(n2804), .A2(\bank_register[8][5] ), .B1(n2801), .B2(
        \bank_register[16][5] ), .ZN(n2046) );
  AOI22_X1 U1087 ( .A1(n2886), .A2(\bank_register[22][5] ), .B1(n2876), .B2(
        \bank_register[30][5] ), .ZN(n2028) );
  AOI22_X1 U1088 ( .A1(n2813), .A2(\bank_register[4][6] ), .B1(n3240), .B2(
        n2014), .ZN(n2013) );
  NAND2_X1 U1089 ( .A1(n2015), .A2(n2016), .ZN(n2014) );
  AOI221_X1 U1090 ( .B1(n2885), .B2(\bank_register[21][6] ), .C1(n2874), .C2(
        \bank_register[29][6] ), .A(n2018), .ZN(n2015) );
  AOI221_X1 U1091 ( .B1(n2841), .B2(\bank_register[25][6] ), .C1(n2830), .C2(
        \bank_register[13][6] ), .A(n2017), .ZN(n2016) );
  AOI22_X1 U1092 ( .A1(n2804), .A2(\bank_register[8][6] ), .B1(n2801), .B2(
        \bank_register[16][6] ), .ZN(n2021) );
  AOI22_X1 U1093 ( .A1(n2887), .A2(\bank_register[22][6] ), .B1(n2875), .B2(
        \bank_register[30][6] ), .ZN(n2003) );
  AOI22_X1 U1094 ( .A1(n2813), .A2(\bank_register[4][7] ), .B1(n3240), .B2(
        n1989), .ZN(n1988) );
  NAND2_X1 U1095 ( .A1(n1990), .A2(n1991), .ZN(n1989) );
  AOI221_X1 U1096 ( .B1(n2884), .B2(\bank_register[21][7] ), .C1(n2873), .C2(
        \bank_register[29][7] ), .A(n1993), .ZN(n1990) );
  AOI221_X1 U1097 ( .B1(n2840), .B2(\bank_register[25][7] ), .C1(n2829), .C2(
        \bank_register[13][7] ), .A(n1992), .ZN(n1991) );
  AOI22_X1 U1098 ( .A1(n2804), .A2(\bank_register[8][7] ), .B1(n2801), .B2(
        \bank_register[16][7] ), .ZN(n1996) );
  AOI22_X1 U1099 ( .A1(n2887), .A2(\bank_register[22][7] ), .B1(n2875), .B2(
        \bank_register[30][7] ), .ZN(n1978) );
  AOI22_X1 U1100 ( .A1(n2813), .A2(\bank_register[4][8] ), .B1(
        read_address_1[0]), .B2(n1964), .ZN(n1963) );
  NAND2_X1 U1101 ( .A1(n1965), .A2(n1966), .ZN(n1964) );
  AOI221_X1 U1102 ( .B1(n2884), .B2(\bank_register[21][8] ), .C1(n2873), .C2(
        \bank_register[29][8] ), .A(n1968), .ZN(n1965) );
  AOI221_X1 U1103 ( .B1(n2840), .B2(\bank_register[25][8] ), .C1(n2829), .C2(
        \bank_register[13][8] ), .A(n1967), .ZN(n1966) );
  AOI22_X1 U1104 ( .A1(n2804), .A2(\bank_register[8][8] ), .B1(n2801), .B2(
        \bank_register[16][8] ), .ZN(n1971) );
  AOI22_X1 U1105 ( .A1(n2886), .A2(\bank_register[22][8] ), .B1(n2877), .B2(
        \bank_register[30][8] ), .ZN(n1953) );
  AOI22_X1 U1106 ( .A1(n2813), .A2(\bank_register[4][9] ), .B1(n3240), .B2(
        n1935), .ZN(n1933) );
  NAND2_X1 U1107 ( .A1(n1936), .A2(n1937), .ZN(n1935) );
  AOI221_X1 U1108 ( .B1(n2884), .B2(\bank_register[21][9] ), .C1(n2873), .C2(
        \bank_register[29][9] ), .A(n1939), .ZN(n1936) );
  AOI221_X1 U1109 ( .B1(n2840), .B2(\bank_register[25][9] ), .C1(n2829), .C2(
        \bank_register[13][9] ), .A(n1938), .ZN(n1937) );
  AOI22_X1 U1110 ( .A1(n2804), .A2(\bank_register[8][9] ), .B1(n2801), .B2(
        \bank_register[16][9] ), .ZN(n1944) );
  AOI22_X1 U1111 ( .A1(n2888), .A2(\bank_register[22][9] ), .B1(n2877), .B2(
        \bank_register[30][9] ), .ZN(n1913) );
  AOI22_X1 U1112 ( .A1(n2811), .A2(\bank_register[4][10] ), .B1(n3240), .B2(
        n2752), .ZN(n2751) );
  NAND2_X1 U1113 ( .A1(n2753), .A2(n2754), .ZN(n2752) );
  AOI221_X1 U1114 ( .B1(n2884), .B2(\bank_register[21][10] ), .C1(n2873), .C2(
        \bank_register[29][10] ), .A(n2756), .ZN(n2753) );
  AOI221_X1 U1115 ( .B1(n2840), .B2(\bank_register[25][10] ), .C1(n2829), .C2(
        \bank_register[13][10] ), .A(n2755), .ZN(n2754) );
  AOI22_X1 U1116 ( .A1(n2802), .A2(\bank_register[8][10] ), .B1(n2767), .B2(
        \bank_register[16][10] ), .ZN(n2759) );
  AOI22_X1 U1117 ( .A1(n2891), .A2(\bank_register[22][10] ), .B1(n2880), .B2(
        \bank_register[30][10] ), .ZN(n2741) );
  AOI22_X1 U1118 ( .A1(n2811), .A2(\bank_register[4][11] ), .B1(n3240), .B2(
        n2727), .ZN(n2726) );
  NAND2_X1 U1119 ( .A1(n2728), .A2(n2729), .ZN(n2727) );
  AOI221_X1 U1120 ( .B1(n2884), .B2(\bank_register[21][11] ), .C1(n2873), .C2(
        \bank_register[29][11] ), .A(n2731), .ZN(n2728) );
  AOI221_X1 U1121 ( .B1(n2840), .B2(\bank_register[25][11] ), .C1(n2829), .C2(
        \bank_register[13][11] ), .A(n2730), .ZN(n2729) );
  AOI22_X1 U1122 ( .A1(n2802), .A2(\bank_register[8][11] ), .B1(n2767), .B2(
        \bank_register[16][11] ), .ZN(n2734) );
  AOI22_X1 U1123 ( .A1(n2891), .A2(\bank_register[22][11] ), .B1(n2880), .B2(
        \bank_register[30][11] ), .ZN(n2716) );
  AOI22_X1 U1124 ( .A1(n2811), .A2(\bank_register[4][12] ), .B1(n3240), .B2(
        n2702), .ZN(n2701) );
  NAND2_X1 U1125 ( .A1(n2703), .A2(n2704), .ZN(n2702) );
  AOI221_X1 U1126 ( .B1(n2884), .B2(\bank_register[21][12] ), .C1(n2873), .C2(
        \bank_register[29][12] ), .A(n2706), .ZN(n2703) );
  AOI221_X1 U1127 ( .B1(n2840), .B2(\bank_register[25][12] ), .C1(n2829), .C2(
        \bank_register[13][12] ), .A(n2705), .ZN(n2704) );
  AOI22_X1 U1128 ( .A1(n2802), .A2(\bank_register[8][12] ), .B1(n2767), .B2(
        \bank_register[16][12] ), .ZN(n2709) );
  AOI22_X1 U1129 ( .A1(n2891), .A2(\bank_register[22][12] ), .B1(n2880), .B2(
        \bank_register[30][12] ), .ZN(n2691) );
  AOI22_X1 U1130 ( .A1(n2811), .A2(\bank_register[4][13] ), .B1(n3240), .B2(
        n2677), .ZN(n2676) );
  NAND2_X1 U1131 ( .A1(n2678), .A2(n2679), .ZN(n2677) );
  AOI221_X1 U1132 ( .B1(n2884), .B2(\bank_register[21][13] ), .C1(n2873), .C2(
        \bank_register[29][13] ), .A(n2681), .ZN(n2678) );
  AOI221_X1 U1133 ( .B1(n2840), .B2(\bank_register[25][13] ), .C1(n2829), .C2(
        \bank_register[13][13] ), .A(n2680), .ZN(n2679) );
  AOI22_X1 U1134 ( .A1(n2802), .A2(\bank_register[8][13] ), .B1(n2767), .B2(
        \bank_register[16][13] ), .ZN(n2684) );
  AOI22_X1 U1135 ( .A1(n2891), .A2(\bank_register[22][13] ), .B1(n2880), .B2(
        \bank_register[30][13] ), .ZN(n2666) );
  AOI22_X1 U1136 ( .A1(n2811), .A2(\bank_register[4][14] ), .B1(n3240), .B2(
        n2652), .ZN(n2651) );
  NAND2_X1 U1137 ( .A1(n2653), .A2(n2654), .ZN(n2652) );
  AOI221_X1 U1138 ( .B1(n2884), .B2(\bank_register[21][14] ), .C1(n2873), .C2(
        \bank_register[29][14] ), .A(n2656), .ZN(n2653) );
  AOI221_X1 U1139 ( .B1(n2840), .B2(\bank_register[25][14] ), .C1(n2829), .C2(
        \bank_register[13][14] ), .A(n2655), .ZN(n2654) );
  AOI22_X1 U1140 ( .A1(n2802), .A2(\bank_register[8][14] ), .B1(n2767), .B2(
        \bank_register[16][14] ), .ZN(n2659) );
  AOI22_X1 U1141 ( .A1(n2891), .A2(\bank_register[22][14] ), .B1(n2880), .B2(
        \bank_register[30][14] ), .ZN(n2641) );
  AOI22_X1 U1142 ( .A1(n2811), .A2(\bank_register[4][15] ), .B1(n3240), .B2(
        n2627), .ZN(n2626) );
  NAND2_X1 U1143 ( .A1(n2628), .A2(n2629), .ZN(n2627) );
  AOI221_X1 U1144 ( .B1(n2885), .B2(\bank_register[21][15] ), .C1(n2874), .C2(
        \bank_register[29][15] ), .A(n2631), .ZN(n2628) );
  AOI221_X1 U1145 ( .B1(n2841), .B2(\bank_register[25][15] ), .C1(n2830), .C2(
        \bank_register[13][15] ), .A(n2630), .ZN(n2629) );
  AOI22_X1 U1146 ( .A1(n2802), .A2(\bank_register[8][15] ), .B1(n2767), .B2(
        \bank_register[16][15] ), .ZN(n2634) );
  AOI22_X1 U1147 ( .A1(n2890), .A2(\bank_register[22][15] ), .B1(n2880), .B2(
        \bank_register[30][15] ), .ZN(n2616) );
  AOI22_X1 U1148 ( .A1(n2811), .A2(\bank_register[4][16] ), .B1(n3240), .B2(
        n2602), .ZN(n2601) );
  NAND2_X1 U1149 ( .A1(n2603), .A2(n2604), .ZN(n2602) );
  AOI221_X1 U1150 ( .B1(n2884), .B2(\bank_register[21][16] ), .C1(n2874), .C2(
        \bank_register[29][16] ), .A(n2606), .ZN(n2603) );
  AOI221_X1 U1151 ( .B1(n2840), .B2(\bank_register[25][16] ), .C1(n2830), .C2(
        \bank_register[13][16] ), .A(n2605), .ZN(n2604) );
  AOI22_X1 U1152 ( .A1(n2802), .A2(\bank_register[8][16] ), .B1(n2767), .B2(
        \bank_register[16][16] ), .ZN(n2609) );
  AOI22_X1 U1153 ( .A1(n2890), .A2(\bank_register[22][16] ), .B1(n2879), .B2(
        \bank_register[30][16] ), .ZN(n2591) );
  AOI22_X1 U1154 ( .A1(n2811), .A2(\bank_register[4][17] ), .B1(n3240), .B2(
        n2577), .ZN(n2576) );
  NAND2_X1 U1155 ( .A1(n2578), .A2(n2579), .ZN(n2577) );
  AOI221_X1 U1156 ( .B1(n2885), .B2(\bank_register[21][17] ), .C1(n2873), .C2(
        \bank_register[29][17] ), .A(n2581), .ZN(n2578) );
  AOI221_X1 U1157 ( .B1(n2841), .B2(\bank_register[25][17] ), .C1(n2829), .C2(
        \bank_register[13][17] ), .A(n2580), .ZN(n2579) );
  AOI22_X1 U1158 ( .A1(n2802), .A2(\bank_register[8][17] ), .B1(n2767), .B2(
        \bank_register[16][17] ), .ZN(n2584) );
  AOI22_X1 U1159 ( .A1(n2890), .A2(\bank_register[22][17] ), .B1(n2879), .B2(
        \bank_register[30][17] ), .ZN(n2566) );
  AOI22_X1 U1160 ( .A1(n2811), .A2(\bank_register[4][18] ), .B1(n3240), .B2(
        n2552), .ZN(n2551) );
  NAND2_X1 U1161 ( .A1(n2553), .A2(n2554), .ZN(n2552) );
  AOI221_X1 U1162 ( .B1(n2885), .B2(\bank_register[21][18] ), .C1(n2874), .C2(
        \bank_register[29][18] ), .A(n2556), .ZN(n2553) );
  AOI221_X1 U1163 ( .B1(n2841), .B2(\bank_register[25][18] ), .C1(n2830), .C2(
        \bank_register[13][18] ), .A(n2555), .ZN(n2554) );
  AOI22_X1 U1164 ( .A1(n2802), .A2(\bank_register[8][18] ), .B1(n2767), .B2(
        \bank_register[16][18] ), .ZN(n2559) );
  AOI22_X1 U1165 ( .A1(n2890), .A2(\bank_register[22][18] ), .B1(n2879), .B2(
        \bank_register[30][18] ), .ZN(n2541) );
  AOI22_X1 U1166 ( .A1(n2811), .A2(\bank_register[4][19] ), .B1(
        read_address_1[0]), .B2(n2527), .ZN(n2526) );
  NAND2_X1 U1167 ( .A1(n2528), .A2(n2529), .ZN(n2527) );
  AOI221_X1 U1168 ( .B1(n2885), .B2(\bank_register[21][19] ), .C1(n2875), .C2(
        \bank_register[29][19] ), .A(n2531), .ZN(n2528) );
  AOI221_X1 U1169 ( .B1(n2841), .B2(\bank_register[25][19] ), .C1(n2831), .C2(
        \bank_register[13][19] ), .A(n2530), .ZN(n2529) );
  AOI22_X1 U1170 ( .A1(n2802), .A2(\bank_register[8][19] ), .B1(n2767), .B2(
        \bank_register[16][19] ), .ZN(n2534) );
  AOI22_X1 U1171 ( .A1(n2890), .A2(\bank_register[22][19] ), .B1(n2879), .B2(
        \bank_register[30][19] ), .ZN(n2516) );
  AOI22_X1 U1172 ( .A1(n2812), .A2(\bank_register[4][20] ), .B1(
        read_address_1[0]), .B2(n2477), .ZN(n2476) );
  NAND2_X1 U1173 ( .A1(n2478), .A2(n2479), .ZN(n2477) );
  AOI221_X1 U1174 ( .B1(n2886), .B2(\bank_register[21][20] ), .C1(n2875), .C2(
        \bank_register[29][20] ), .A(n2481), .ZN(n2478) );
  AOI221_X1 U1175 ( .B1(n2842), .B2(\bank_register[25][20] ), .C1(n2831), .C2(
        \bank_register[13][20] ), .A(n2480), .ZN(n2479) );
  AOI22_X1 U1176 ( .A1(n2803), .A2(\bank_register[8][20] ), .B1(n2800), .B2(
        \bank_register[16][20] ), .ZN(n2484) );
  AOI22_X1 U1177 ( .A1(n2889), .A2(\bank_register[22][20] ), .B1(n2879), .B2(
        \bank_register[30][20] ), .ZN(n2466) );
  AOI22_X1 U1178 ( .A1(n2812), .A2(\bank_register[4][21] ), .B1(
        read_address_1[0]), .B2(n2452), .ZN(n2451) );
  NAND2_X1 U1179 ( .A1(n2453), .A2(n2454), .ZN(n2452) );
  AOI221_X1 U1180 ( .B1(n2885), .B2(\bank_register[21][21] ), .C1(n2874), .C2(
        \bank_register[29][21] ), .A(n2456), .ZN(n2453) );
  AOI221_X1 U1181 ( .B1(n2841), .B2(\bank_register[25][21] ), .C1(n2830), .C2(
        \bank_register[13][21] ), .A(n2455), .ZN(n2454) );
  AOI22_X1 U1182 ( .A1(n2803), .A2(\bank_register[8][21] ), .B1(n2800), .B2(
        \bank_register[16][21] ), .ZN(n2459) );
  AOI22_X1 U1183 ( .A1(n2889), .A2(\bank_register[22][21] ), .B1(n2878), .B2(
        \bank_register[30][21] ), .ZN(n2441) );
  AOI22_X1 U1184 ( .A1(n2812), .A2(\bank_register[4][22] ), .B1(
        read_address_1[0]), .B2(n2427), .ZN(n2426) );
  NAND2_X1 U1185 ( .A1(n2428), .A2(n2429), .ZN(n2427) );
  AOI221_X1 U1186 ( .B1(n2886), .B2(\bank_register[21][22] ), .C1(n2874), .C2(
        \bank_register[29][22] ), .A(n2431), .ZN(n2428) );
  AOI221_X1 U1187 ( .B1(n2842), .B2(\bank_register[25][22] ), .C1(n2830), .C2(
        \bank_register[13][22] ), .A(n2430), .ZN(n2429) );
  AOI22_X1 U1188 ( .A1(n2803), .A2(\bank_register[8][22] ), .B1(n2800), .B2(
        \bank_register[16][22] ), .ZN(n2434) );
  AOI22_X1 U1189 ( .A1(n2889), .A2(\bank_register[22][22] ), .B1(n2878), .B2(
        \bank_register[30][22] ), .ZN(n2416) );
  AOI22_X1 U1190 ( .A1(n2812), .A2(\bank_register[4][23] ), .B1(
        read_address_1[0]), .B2(n2402), .ZN(n2401) );
  NAND2_X1 U1191 ( .A1(n2403), .A2(n2404), .ZN(n2402) );
  AOI221_X1 U1192 ( .B1(n2885), .B2(\bank_register[21][23] ), .C1(n2874), .C2(
        \bank_register[29][23] ), .A(n2406), .ZN(n2403) );
  AOI221_X1 U1193 ( .B1(n2841), .B2(\bank_register[25][23] ), .C1(n2830), .C2(
        \bank_register[13][23] ), .A(n2405), .ZN(n2404) );
  AOI22_X1 U1194 ( .A1(n2803), .A2(\bank_register[8][23] ), .B1(n2800), .B2(
        \bank_register[16][23] ), .ZN(n2409) );
  AOI22_X1 U1195 ( .A1(n2889), .A2(\bank_register[22][23] ), .B1(n2878), .B2(
        \bank_register[30][23] ), .ZN(n2391) );
  AOI22_X1 U1196 ( .A1(n2812), .A2(\bank_register[4][24] ), .B1(
        read_address_1[0]), .B2(n2377), .ZN(n2376) );
  NAND2_X1 U1197 ( .A1(n2378), .A2(n2379), .ZN(n2377) );
  AOI221_X1 U1198 ( .B1(n2886), .B2(\bank_register[21][24] ), .C1(n2875), .C2(
        \bank_register[29][24] ), .A(n2381), .ZN(n2378) );
  AOI221_X1 U1199 ( .B1(n2842), .B2(\bank_register[25][24] ), .C1(n2831), .C2(
        \bank_register[13][24] ), .A(n2380), .ZN(n2379) );
  AOI22_X1 U1200 ( .A1(n2803), .A2(\bank_register[8][24] ), .B1(n2800), .B2(
        \bank_register[16][24] ), .ZN(n2384) );
  AOI22_X1 U1201 ( .A1(n2889), .A2(\bank_register[22][24] ), .B1(n2878), .B2(
        \bank_register[30][24] ), .ZN(n2364) );
  AOI22_X1 U1202 ( .A1(n2812), .A2(\bank_register[4][25] ), .B1(
        read_address_1[0]), .B2(n2346), .ZN(n2344) );
  NAND2_X1 U1203 ( .A1(n2347), .A2(n2348), .ZN(n2346) );
  AOI221_X1 U1204 ( .B1(n2885), .B2(\bank_register[21][25] ), .C1(n2875), .C2(
        \bank_register[29][25] ), .A(n2351), .ZN(n2347) );
  AOI221_X1 U1205 ( .B1(n2841), .B2(\bank_register[25][25] ), .C1(n2831), .C2(
        \bank_register[13][25] ), .A(n2350), .ZN(n2348) );
  AOI22_X1 U1206 ( .A1(n2803), .A2(\bank_register[8][25] ), .B1(n2800), .B2(
        \bank_register[16][25] ), .ZN(n2355) );
  AOI22_X1 U1207 ( .A1(n2889), .A2(\bank_register[22][25] ), .B1(n2878), .B2(
        \bank_register[30][25] ), .ZN(n2331) );
  AOI22_X1 U1208 ( .A1(n2812), .A2(\bank_register[4][26] ), .B1(
        read_address_1[0]), .B2(n2312), .ZN(n2311) );
  NAND2_X1 U1209 ( .A1(n2314), .A2(n2315), .ZN(n2312) );
  AOI221_X1 U1210 ( .B1(n2886), .B2(\bank_register[21][26] ), .C1(n2875), .C2(
        \bank_register[29][26] ), .A(n2318), .ZN(n2314) );
  AOI221_X1 U1211 ( .B1(n2842), .B2(\bank_register[25][26] ), .C1(n2831), .C2(
        \bank_register[13][26] ), .A(n2316), .ZN(n2315) );
  AOI22_X1 U1212 ( .A1(n2803), .A2(\bank_register[8][26] ), .B1(n2800), .B2(
        \bank_register[16][26] ), .ZN(n2322) );
  AOI22_X1 U1213 ( .A1(n2888), .A2(\bank_register[22][26] ), .B1(n2878), .B2(
        \bank_register[30][26] ), .ZN(n2298) );
  AOI22_X1 U1214 ( .A1(n2812), .A2(\bank_register[4][27] ), .B1(
        read_address_1[0]), .B2(n2279), .ZN(n2278) );
  NAND2_X1 U1215 ( .A1(n2280), .A2(n2282), .ZN(n2279) );
  AOI221_X1 U1216 ( .B1(n2885), .B2(\bank_register[21][27] ), .C1(n2874), .C2(
        \bank_register[29][27] ), .A(n2284), .ZN(n2280) );
  AOI221_X1 U1217 ( .B1(n2841), .B2(\bank_register[25][27] ), .C1(n2830), .C2(
        \bank_register[13][27] ), .A(n2283), .ZN(n2282) );
  AOI22_X1 U1218 ( .A1(n2803), .A2(\bank_register[8][27] ), .B1(n2800), .B2(
        \bank_register[16][27] ), .ZN(n2288) );
  AOI22_X1 U1219 ( .A1(n2888), .A2(\bank_register[22][27] ), .B1(n2877), .B2(
        \bank_register[30][27] ), .ZN(n2264) );
  AOI22_X1 U1220 ( .A1(n2812), .A2(\bank_register[4][28] ), .B1(
        read_address_1[0]), .B2(n2246), .ZN(n2244) );
  NAND2_X1 U1221 ( .A1(n2247), .A2(n2248), .ZN(n2246) );
  AOI221_X1 U1222 ( .B1(n2886), .B2(\bank_register[21][28] ), .C1(n2875), .C2(
        \bank_register[29][28] ), .A(n2251), .ZN(n2247) );
  AOI221_X1 U1223 ( .B1(n2842), .B2(\bank_register[25][28] ), .C1(n2831), .C2(
        \bank_register[13][28] ), .A(n2250), .ZN(n2248) );
  AOI22_X1 U1224 ( .A1(n2803), .A2(\bank_register[8][28] ), .B1(n2800), .B2(
        \bank_register[16][28] ), .ZN(n2255) );
  AOI22_X1 U1225 ( .A1(n2888), .A2(\bank_register[22][28] ), .B1(n2877), .B2(
        \bank_register[30][28] ), .ZN(n2229) );
  AOI22_X1 U1226 ( .A1(n2812), .A2(\bank_register[4][29] ), .B1(
        read_address_1[0]), .B2(n2208), .ZN(n2207) );
  NAND2_X1 U1227 ( .A1(n2210), .A2(n2211), .ZN(n2208) );
  AOI221_X1 U1228 ( .B1(n2886), .B2(\bank_register[21][29] ), .C1(n2874), .C2(
        \bank_register[29][29] ), .A(n2214), .ZN(n2210) );
  AOI221_X1 U1229 ( .B1(n2842), .B2(\bank_register[25][29] ), .C1(n2830), .C2(
        \bank_register[13][29] ), .A(n2213), .ZN(n2211) );
  AOI22_X1 U1230 ( .A1(n2803), .A2(\bank_register[8][29] ), .B1(n2800), .B2(
        \bank_register[16][29] ), .ZN(n2219) );
  AOI22_X1 U1231 ( .A1(n2888), .A2(\bank_register[22][29] ), .B1(n2877), .B2(
        \bank_register[30][29] ), .ZN(n2192) );
  AOI22_X1 U1232 ( .A1(n2812), .A2(\bank_register[4][30] ), .B1(
        read_address_1[0]), .B2(n2139), .ZN(n2138) );
  NAND2_X1 U1233 ( .A1(n2140), .A2(n2141), .ZN(n2139) );
  AOI221_X1 U1234 ( .B1(n2885), .B2(\bank_register[21][30] ), .C1(n2875), .C2(
        \bank_register[29][30] ), .A(n2143), .ZN(n2140) );
  AOI221_X1 U1235 ( .B1(n2841), .B2(\bank_register[25][30] ), .C1(n2831), .C2(
        \bank_register[13][30] ), .A(n2142), .ZN(n2141) );
  AOI22_X1 U1236 ( .A1(n2803), .A2(\bank_register[8][30] ), .B1(n2800), .B2(
        \bank_register[16][30] ), .ZN(n2146) );
  AOI22_X1 U1237 ( .A1(n2887), .A2(\bank_register[22][30] ), .B1(n2876), .B2(
        \bank_register[30][30] ), .ZN(n2128) );
  AOI22_X1 U1238 ( .A1(n2813), .A2(\bank_register[4][31] ), .B1(
        read_address_1[0]), .B2(n2114), .ZN(n2113) );
  NAND2_X1 U1239 ( .A1(n2115), .A2(n2116), .ZN(n2114) );
  AOI221_X1 U1240 ( .B1(n2886), .B2(\bank_register[21][31] ), .C1(n2874), .C2(
        \bank_register[29][31] ), .A(n2118), .ZN(n2115) );
  AOI221_X1 U1241 ( .B1(n2842), .B2(\bank_register[25][31] ), .C1(n2830), .C2(
        \bank_register[13][31] ), .A(n2117), .ZN(n2116) );
  AOI22_X1 U1242 ( .A1(n2804), .A2(\bank_register[8][31] ), .B1(n2801), .B2(
        \bank_register[16][31] ), .ZN(n2121) );
  AOI22_X1 U1243 ( .A1(n2887), .A2(\bank_register[22][31] ), .B1(n2877), .B2(
        \bank_register[30][31] ), .ZN(n2103) );
  OAI221_X1 U1244 ( .B1(n1877), .B2(n2865), .C1(n1876), .C2(n2854), .A(n2774), 
        .ZN(n2770) );
  AOI22_X1 U1245 ( .A1(n2847), .A2(\bank_register[27][0] ), .B1(n2832), .B2(
        \bank_register[15][0] ), .ZN(n2774) );
  OAI221_X1 U1246 ( .B1(n1461), .B2(n2911), .C1(n1460), .C2(n2901), .A(n2495), 
        .ZN(n2494) );
  AOI22_X1 U1247 ( .A1(n2890), .A2(\bank_register[23][1] ), .B1(n2879), .B2(
        \bank_register[31][1] ), .ZN(n2495) );
  OAI221_X1 U1248 ( .B1(n1465), .B2(n2868), .C1(n1464), .C2(n2857), .A(n2496), 
        .ZN(n2493) );
  AOI22_X1 U1249 ( .A1(n2846), .A2(\bank_register[27][1] ), .B1(n2835), .B2(
        \bank_register[15][1] ), .ZN(n2496) );
  OAI221_X1 U1250 ( .B1(n1058), .B2(n2866), .C1(n1057), .C2(n2855), .A(n2162), 
        .ZN(n2157) );
  AOI22_X1 U1251 ( .A1(n2844), .A2(\bank_register[27][2] ), .B1(n2833), .B2(
        \bank_register[15][2] ), .ZN(n2162) );
  OAI221_X1 U1252 ( .B1(n947), .B2(n2865), .C1(n946), .C2(n2854), .A(n2083), 
        .ZN(n2080) );
  AOI22_X1 U1253 ( .A1(n2843), .A2(\bank_register[27][3] ), .B1(n2832), .B2(
        \bank_register[15][3] ), .ZN(n2083) );
  OAI221_X1 U1254 ( .B1(n910), .B2(n2865), .C1(n909), .C2(n2854), .A(n2058), 
        .ZN(n2055) );
  AOI22_X1 U1255 ( .A1(n2844), .A2(\bank_register[27][4] ), .B1(n2832), .B2(
        \bank_register[15][4] ), .ZN(n2058) );
  OAI221_X1 U1256 ( .B1(n873), .B2(n2865), .C1(n872), .C2(n2854), .A(n2033), 
        .ZN(n2030) );
  AOI22_X1 U1257 ( .A1(n2843), .A2(\bank_register[27][5] ), .B1(n2832), .B2(
        \bank_register[15][5] ), .ZN(n2033) );
  OAI221_X1 U1258 ( .B1(n799), .B2(n2865), .C1(n798), .C2(n2854), .A(n1983), 
        .ZN(n1980) );
  AOI22_X1 U1259 ( .A1(n2842), .A2(\bank_register[27][7] ), .B1(n2832), .B2(
        \bank_register[15][7] ), .ZN(n1983) );
  OAI221_X1 U1260 ( .B1(n762), .B2(n2865), .C1(n761), .C2(n2854), .A(n1958), 
        .ZN(n1955) );
  AOI22_X1 U1261 ( .A1(n2842), .A2(\bank_register[27][8] ), .B1(n2832), .B2(
        \bank_register[15][8] ), .ZN(n1958) );
  OAI221_X1 U1262 ( .B1(n725), .B2(n2865), .C1(n724), .C2(n2855), .A(n1925), 
        .ZN(n1921) );
  AOI22_X1 U1263 ( .A1(n2843), .A2(\bank_register[27][9] ), .B1(n2833), .B2(
        \bank_register[15][9] ), .ZN(n1925) );
  OAI221_X1 U1264 ( .B1(n1831), .B2(n2913), .C1(n1830), .C2(n2902), .A(n2745), 
        .ZN(n2744) );
  AOI22_X1 U1265 ( .A1(n2891), .A2(\bank_register[23][10] ), .B1(n2880), .B2(
        \bank_register[31][10] ), .ZN(n2745) );
  OAI221_X1 U1266 ( .B1(n1835), .B2(n2869), .C1(n1834), .C2(n2858), .A(n2746), 
        .ZN(n2743) );
  AOI22_X1 U1267 ( .A1(n2847), .A2(\bank_register[27][10] ), .B1(n2836), .B2(
        \bank_register[15][10] ), .ZN(n2746) );
  OAI221_X1 U1268 ( .B1(n1794), .B2(n2913), .C1(n1793), .C2(n2902), .A(n2720), 
        .ZN(n2719) );
  AOI22_X1 U1269 ( .A1(n2891), .A2(\bank_register[23][11] ), .B1(n2880), .B2(
        \bank_register[31][11] ), .ZN(n2720) );
  OAI221_X1 U1270 ( .B1(n1798), .B2(n2869), .C1(n1797), .C2(n2858), .A(n2721), 
        .ZN(n2718) );
  AOI22_X1 U1271 ( .A1(n2847), .A2(\bank_register[27][11] ), .B1(n2836), .B2(
        \bank_register[15][11] ), .ZN(n2721) );
  OAI221_X1 U1272 ( .B1(n1757), .B2(n2913), .C1(n1756), .C2(n2902), .A(n2695), 
        .ZN(n2694) );
  AOI22_X1 U1273 ( .A1(n2891), .A2(\bank_register[23][12] ), .B1(n2880), .B2(
        \bank_register[31][12] ), .ZN(n2695) );
  OAI221_X1 U1274 ( .B1(n1761), .B2(n2869), .C1(n1760), .C2(n2858), .A(n2696), 
        .ZN(n2693) );
  AOI22_X1 U1275 ( .A1(n2847), .A2(\bank_register[27][12] ), .B1(n2836), .B2(
        \bank_register[15][12] ), .ZN(n2696) );
  OAI221_X1 U1276 ( .B1(n1720), .B2(n2913), .C1(n1719), .C2(n2902), .A(n2670), 
        .ZN(n2669) );
  AOI22_X1 U1277 ( .A1(n2891), .A2(\bank_register[23][13] ), .B1(n2880), .B2(
        \bank_register[31][13] ), .ZN(n2670) );
  OAI221_X1 U1278 ( .B1(n1724), .B2(n2869), .C1(n1723), .C2(n2858), .A(n2671), 
        .ZN(n2668) );
  AOI22_X1 U1279 ( .A1(n2847), .A2(\bank_register[27][13] ), .B1(n2836), .B2(
        \bank_register[15][13] ), .ZN(n2671) );
  OAI221_X1 U1280 ( .B1(n1683), .B2(n2912), .C1(n1682), .C2(n2902), .A(n2645), 
        .ZN(n2644) );
  AOI22_X1 U1281 ( .A1(n2891), .A2(\bank_register[23][14] ), .B1(n2880), .B2(
        \bank_register[31][14] ), .ZN(n2645) );
  OAI221_X1 U1282 ( .B1(n1687), .B2(n2868), .C1(n1686), .C2(n2858), .A(n2646), 
        .ZN(n2643) );
  AOI22_X1 U1283 ( .A1(n2847), .A2(\bank_register[27][14] ), .B1(n2836), .B2(
        \bank_register[15][14] ), .ZN(n2646) );
  OAI221_X1 U1284 ( .B1(n1646), .B2(n2912), .C1(n1645), .C2(n2902), .A(n2620), 
        .ZN(n2619) );
  AOI22_X1 U1285 ( .A1(n2890), .A2(\bank_register[23][15] ), .B1(n2880), .B2(
        \bank_register[31][15] ), .ZN(n2620) );
  OAI221_X1 U1286 ( .B1(n1650), .B2(n2868), .C1(n1649), .C2(n2858), .A(n2621), 
        .ZN(n2618) );
  AOI22_X1 U1287 ( .A1(n2846), .A2(\bank_register[27][15] ), .B1(n2836), .B2(
        \bank_register[15][15] ), .ZN(n2621) );
  OAI221_X1 U1288 ( .B1(n1609), .B2(n2912), .C1(n1608), .C2(n2901), .A(n2595), 
        .ZN(n2594) );
  AOI22_X1 U1289 ( .A1(n2890), .A2(\bank_register[23][16] ), .B1(n2879), .B2(
        \bank_register[31][16] ), .ZN(n2595) );
  OAI221_X1 U1290 ( .B1(n1613), .B2(n2868), .C1(n1612), .C2(n2857), .A(n2596), 
        .ZN(n2593) );
  AOI22_X1 U1291 ( .A1(n2846), .A2(\bank_register[27][16] ), .B1(n2835), .B2(
        \bank_register[15][16] ), .ZN(n2596) );
  OAI221_X1 U1292 ( .B1(n1572), .B2(n2912), .C1(n1571), .C2(n2901), .A(n2570), 
        .ZN(n2569) );
  AOI22_X1 U1293 ( .A1(n2890), .A2(\bank_register[23][17] ), .B1(n2879), .B2(
        \bank_register[31][17] ), .ZN(n2570) );
  OAI221_X1 U1294 ( .B1(n1576), .B2(n2868), .C1(n1575), .C2(n2857), .A(n2571), 
        .ZN(n2568) );
  AOI22_X1 U1295 ( .A1(n2846), .A2(\bank_register[27][17] ), .B1(n2835), .B2(
        \bank_register[15][17] ), .ZN(n2571) );
  OAI221_X1 U1296 ( .B1(n1535), .B2(n2912), .C1(n1534), .C2(n2901), .A(n2545), 
        .ZN(n2544) );
  AOI22_X1 U1297 ( .A1(n2890), .A2(\bank_register[23][18] ), .B1(n2879), .B2(
        \bank_register[31][18] ), .ZN(n2545) );
  OAI221_X1 U1298 ( .B1(n1539), .B2(n2868), .C1(n1538), .C2(n2857), .A(n2546), 
        .ZN(n2543) );
  AOI22_X1 U1299 ( .A1(n2846), .A2(\bank_register[27][18] ), .B1(n2835), .B2(
        \bank_register[15][18] ), .ZN(n2546) );
  OAI221_X1 U1300 ( .B1(n1498), .B2(n2912), .C1(n1497), .C2(n2901), .A(n2520), 
        .ZN(n2519) );
  AOI22_X1 U1301 ( .A1(n2890), .A2(\bank_register[23][19] ), .B1(n2879), .B2(
        \bank_register[31][19] ), .ZN(n2520) );
  OAI221_X1 U1302 ( .B1(n1502), .B2(n2868), .C1(n1501), .C2(n2857), .A(n2521), 
        .ZN(n2518) );
  AOI22_X1 U1303 ( .A1(n2846), .A2(\bank_register[27][19] ), .B1(n2835), .B2(
        \bank_register[15][19] ), .ZN(n2521) );
  OAI221_X1 U1304 ( .B1(n1424), .B2(n2911), .C1(n1423), .C2(n2901), .A(n2470), 
        .ZN(n2469) );
  AOI22_X1 U1305 ( .A1(n2889), .A2(\bank_register[23][20] ), .B1(n2879), .B2(
        \bank_register[31][20] ), .ZN(n2470) );
  OAI221_X1 U1306 ( .B1(n1391), .B2(n2867), .C1(n1390), .C2(n2856), .A(n2446), 
        .ZN(n2443) );
  AOI22_X1 U1307 ( .A1(n2845), .A2(\bank_register[27][21] ), .B1(n2834), .B2(
        \bank_register[15][21] ), .ZN(n2446) );
  OAI221_X1 U1308 ( .B1(n1354), .B2(n2867), .C1(n1353), .C2(n2856), .A(n2421), 
        .ZN(n2418) );
  AOI22_X1 U1309 ( .A1(n2845), .A2(\bank_register[27][22] ), .B1(n2834), .B2(
        \bank_register[15][22] ), .ZN(n2421) );
  OAI221_X1 U1310 ( .B1(n1317), .B2(n2867), .C1(n1316), .C2(n2856), .A(n2396), 
        .ZN(n2393) );
  AOI22_X1 U1311 ( .A1(n2845), .A2(\bank_register[27][23] ), .B1(n2834), .B2(
        \bank_register[15][23] ), .ZN(n2396) );
  OAI221_X1 U1312 ( .B1(n1280), .B2(n2867), .C1(n1279), .C2(n2856), .A(n2371), 
        .ZN(n2367) );
  AOI22_X1 U1313 ( .A1(n2845), .A2(\bank_register[27][24] ), .B1(n2834), .B2(
        \bank_register[15][24] ), .ZN(n2371) );
  OAI221_X1 U1314 ( .B1(n1243), .B2(n2867), .C1(n1242), .C2(n2856), .A(n2338), 
        .ZN(n2334) );
  AOI22_X1 U1315 ( .A1(n2845), .A2(\bank_register[27][25] ), .B1(n2834), .B2(
        \bank_register[15][25] ), .ZN(n2338) );
  OAI221_X1 U1316 ( .B1(n1206), .B2(n2866), .C1(n1205), .C2(n2856), .A(n2304), 
        .ZN(n2300) );
  AOI22_X1 U1317 ( .A1(n2844), .A2(\bank_register[27][26] ), .B1(n2834), .B2(
        \bank_register[15][26] ), .ZN(n2304) );
  OAI221_X1 U1318 ( .B1(n1169), .B2(n2866), .C1(n1168), .C2(n2855), .A(n2271), 
        .ZN(n2267) );
  AOI22_X1 U1319 ( .A1(n2844), .A2(\bank_register[27][27] ), .B1(n2833), .B2(
        \bank_register[15][27] ), .ZN(n2271) );
  OAI221_X1 U1320 ( .B1(n1132), .B2(n2866), .C1(n1131), .C2(n2855), .A(n2237), 
        .ZN(n2232) );
  AOI22_X1 U1321 ( .A1(n2844), .A2(\bank_register[27][28] ), .B1(n2833), .B2(
        \bank_register[15][28] ), .ZN(n2237) );
  OAI221_X1 U1322 ( .B1(n1095), .B2(n2866), .C1(n1094), .C2(n2855), .A(n2199), 
        .ZN(n2195) );
  AOI22_X1 U1323 ( .A1(n2844), .A2(\bank_register[27][29] ), .B1(n2833), .B2(
        \bank_register[15][29] ), .ZN(n2199) );
  OAI221_X1 U1324 ( .B1(n1021), .B2(n2865), .C1(n1020), .C2(n2854), .A(n2133), 
        .ZN(n2130) );
  AOI22_X1 U1325 ( .A1(n2844), .A2(\bank_register[27][30] ), .B1(n2832), .B2(
        \bank_register[15][30] ), .ZN(n2133) );
  OAI221_X1 U1326 ( .B1(n984), .B2(n2865), .C1(n983), .C2(n2854), .A(n2108), 
        .ZN(n2105) );
  AOI22_X1 U1327 ( .A1(n2843), .A2(\bank_register[27][31] ), .B1(n2832), .B2(
        \bank_register[15][31] ), .ZN(n2108) );
  AOI22_X1 U1328 ( .A1(\bank_register[4][0] ), .A2(n3009), .B1(
        read_address_2[0]), .B2(n1858), .ZN(n1850) );
  NAND2_X1 U1329 ( .A1(n1859), .A2(n1860), .ZN(n1858) );
  AOI221_X1 U1330 ( .B1(\bank_register[21][0] ), .B2(n2958), .C1(
        \bank_register[29][0] ), .C2(n2947), .A(n1864), .ZN(n1859) );
  AOI221_X1 U1331 ( .B1(\bank_register[25][0] ), .B2(n3002), .C1(
        \bank_register[13][0] ), .C2(n2991), .A(n1861), .ZN(n1860) );
  AOI22_X1 U1332 ( .A1(\bank_register[4][10] ), .A2(n3009), .B1(n3238), .B2(
        n1817), .ZN(n1813) );
  NAND2_X1 U1333 ( .A1(n1818), .A2(n1819), .ZN(n1817) );
  AOI221_X1 U1334 ( .B1(\bank_register[21][10] ), .B2(n2958), .C1(
        \bank_register[29][10] ), .C2(n2947), .A(n1823), .ZN(n1818) );
  AOI221_X1 U1335 ( .B1(\bank_register[25][10] ), .B2(n3002), .C1(
        \bank_register[13][10] ), .C2(n2991), .A(n1820), .ZN(n1819) );
  AOI22_X1 U1336 ( .A1(\bank_register[4][11] ), .A2(n3009), .B1(n3238), .B2(
        n1780), .ZN(n1776) );
  NAND2_X1 U1337 ( .A1(n1781), .A2(n1782), .ZN(n1780) );
  AOI221_X1 U1338 ( .B1(\bank_register[21][11] ), .B2(n2958), .C1(
        \bank_register[29][11] ), .C2(n2947), .A(n1786), .ZN(n1781) );
  AOI221_X1 U1339 ( .B1(\bank_register[25][11] ), .B2(n3002), .C1(
        \bank_register[13][11] ), .C2(n2991), .A(n1783), .ZN(n1782) );
  AOI22_X1 U1340 ( .A1(\bank_register[4][12] ), .A2(n3009), .B1(n3238), .B2(
        n1743), .ZN(n1739) );
  NAND2_X1 U1341 ( .A1(n1744), .A2(n1745), .ZN(n1743) );
  AOI221_X1 U1342 ( .B1(\bank_register[21][12] ), .B2(n2958), .C1(
        \bank_register[29][12] ), .C2(n2947), .A(n1749), .ZN(n1744) );
  AOI221_X1 U1343 ( .B1(\bank_register[25][12] ), .B2(n3002), .C1(
        \bank_register[13][12] ), .C2(n2991), .A(n1746), .ZN(n1745) );
  AOI22_X1 U1344 ( .A1(\bank_register[4][13] ), .A2(n3009), .B1(n3238), .B2(
        n1706), .ZN(n1702) );
  NAND2_X1 U1345 ( .A1(n1707), .A2(n1708), .ZN(n1706) );
  AOI221_X1 U1346 ( .B1(\bank_register[21][13] ), .B2(n2958), .C1(
        \bank_register[29][13] ), .C2(n2947), .A(n1712), .ZN(n1707) );
  AOI221_X1 U1347 ( .B1(\bank_register[25][13] ), .B2(n3002), .C1(
        \bank_register[13][13] ), .C2(n2991), .A(n1709), .ZN(n1708) );
  AOI22_X1 U1348 ( .A1(\bank_register[4][14] ), .A2(n3009), .B1(n3238), .B2(
        n1669), .ZN(n1665) );
  NAND2_X1 U1349 ( .A1(n1670), .A2(n1671), .ZN(n1669) );
  AOI221_X1 U1350 ( .B1(\bank_register[21][14] ), .B2(n2958), .C1(
        \bank_register[29][14] ), .C2(n2947), .A(n1675), .ZN(n1670) );
  AOI221_X1 U1351 ( .B1(\bank_register[25][14] ), .B2(n3002), .C1(
        \bank_register[13][14] ), .C2(n2991), .A(n1672), .ZN(n1671) );
  AOI22_X1 U1352 ( .A1(\bank_register[4][15] ), .A2(n3009), .B1(n3238), .B2(
        n1632), .ZN(n1628) );
  NAND2_X1 U1353 ( .A1(n1633), .A2(n1634), .ZN(n1632) );
  AOI221_X1 U1354 ( .B1(\bank_register[21][15] ), .B2(n2958), .C1(
        \bank_register[29][15] ), .C2(n2947), .A(n1638), .ZN(n1633) );
  AOI221_X1 U1355 ( .B1(\bank_register[25][15] ), .B2(n3002), .C1(
        \bank_register[13][15] ), .C2(n2991), .A(n1635), .ZN(n1634) );
  AOI22_X1 U1356 ( .A1(\bank_register[4][16] ), .A2(n3009), .B1(n3238), .B2(
        n1595), .ZN(n1591) );
  NAND2_X1 U1357 ( .A1(n1596), .A2(n1597), .ZN(n1595) );
  AOI221_X1 U1358 ( .B1(\bank_register[21][16] ), .B2(n2958), .C1(
        \bank_register[29][16] ), .C2(n2947), .A(n1601), .ZN(n1596) );
  AOI221_X1 U1359 ( .B1(\bank_register[25][16] ), .B2(n3002), .C1(
        \bank_register[13][16] ), .C2(n2991), .A(n1598), .ZN(n1597) );
  NOR2_X1 U1360 ( .A1(n1888), .A2(read_address_2[4]), .ZN(n1901) );
  NOR2_X1 U1361 ( .A1(n1895), .A2(read_address_2[3]), .ZN(n1898) );
  INV_X1 U1362 ( .A(read_address_2[0]), .ZN(n3239) );
  NOR2_X1 U1363 ( .A1(n2785), .A2(read_address_1[4]), .ZN(n2793) );
  INV_X1 U1364 ( .A(read_address_2[2]), .ZN(n1896) );
  NOR2_X1 U1365 ( .A1(n2786), .A2(read_address_1[3]), .ZN(n2789) );
  NOR2_X1 U1366 ( .A1(n2917), .A2(read_address_1[1]), .ZN(n1928) );
  INV_X1 U1367 ( .A(read_address_1[4]), .ZN(n2786) );
  OAI21_X1 U1368 ( .B1(n2739), .B2(n2740), .A(n2914), .ZN(n2738) );
  OAI221_X1 U1369 ( .B1(n1845), .B2(n2869), .C1(n1844), .C2(n2858), .A(n2742), 
        .ZN(n2739) );
  OAI221_X1 U1370 ( .B1(n1841), .B2(n2913), .C1(n1840), .C2(n2902), .A(n2741), 
        .ZN(n2740) );
  AOI22_X1 U1371 ( .A1(n2847), .A2(\bank_register[26][10] ), .B1(n2836), .B2(
        \bank_register[14][10] ), .ZN(n2742) );
  OAI21_X1 U1372 ( .B1(n2714), .B2(n2715), .A(n2914), .ZN(n2713) );
  OAI221_X1 U1373 ( .B1(n1808), .B2(n2869), .C1(n1807), .C2(n2858), .A(n2717), 
        .ZN(n2714) );
  OAI221_X1 U1374 ( .B1(n1804), .B2(n2913), .C1(n1803), .C2(n2902), .A(n2716), 
        .ZN(n2715) );
  AOI22_X1 U1375 ( .A1(n2847), .A2(\bank_register[26][11] ), .B1(n2836), .B2(
        \bank_register[14][11] ), .ZN(n2717) );
  OAI21_X1 U1376 ( .B1(n2689), .B2(n2690), .A(n2914), .ZN(n2688) );
  OAI221_X1 U1377 ( .B1(n1771), .B2(n2869), .C1(n1770), .C2(n2858), .A(n2692), 
        .ZN(n2689) );
  OAI221_X1 U1378 ( .B1(n1767), .B2(n2913), .C1(n1766), .C2(n2902), .A(n2691), 
        .ZN(n2690) );
  AOI22_X1 U1379 ( .A1(n2847), .A2(\bank_register[26][12] ), .B1(n2836), .B2(
        \bank_register[14][12] ), .ZN(n2692) );
  OAI21_X1 U1380 ( .B1(n2001), .B2(n2002), .A(n2916), .ZN(n2000) );
  OAI221_X1 U1381 ( .B1(n846), .B2(n2864), .C1(n845), .C2(n2853), .A(n2004), 
        .ZN(n2001) );
  OAI221_X1 U1382 ( .B1(n842), .B2(n2908), .C1(n841), .C2(n2897), .A(n2003), 
        .ZN(n2002) );
  AOI22_X1 U1383 ( .A1(n2843), .A2(\bank_register[26][6] ), .B1(n2831), .B2(
        \bank_register[14][6] ), .ZN(n2004) );
  OAI21_X1 U1384 ( .B1(n1976), .B2(n1977), .A(n2916), .ZN(n1975) );
  OAI221_X1 U1385 ( .B1(n809), .B2(n2864), .C1(n808), .C2(n2853), .A(n1979), 
        .ZN(n1976) );
  OAI221_X1 U1386 ( .B1(n805), .B2(n2908), .C1(n804), .C2(n2897), .A(n1978), 
        .ZN(n1977) );
  AOI22_X1 U1387 ( .A1(n2843), .A2(\bank_register[26][7] ), .B1(n2831), .B2(
        \bank_register[14][7] ), .ZN(n1979) );
  OAI21_X1 U1388 ( .B1(n2151), .B2(n2153), .A(n2915), .ZN(n2150) );
  OAI221_X1 U1389 ( .B1(n1068), .B2(n2866), .C1(n1067), .C2(n2855), .A(n2156), 
        .ZN(n2151) );
  OAI221_X1 U1390 ( .B1(n1064), .B2(n2910), .C1(n1063), .C2(n2899), .A(n2154), 
        .ZN(n2153) );
  AOI22_X1 U1391 ( .A1(n2843), .A2(\bank_register[26][2] ), .B1(n2833), .B2(
        \bank_register[14][2] ), .ZN(n2156) );
  OAI21_X1 U1392 ( .B1(n2076), .B2(n2077), .A(n2916), .ZN(n2075) );
  OAI221_X1 U1393 ( .B1(n957), .B2(n2865), .C1(n956), .C2(n2854), .A(n2079), 
        .ZN(n2076) );
  OAI221_X1 U1394 ( .B1(n953), .B2(n2909), .C1(n952), .C2(n2898), .A(n2078), 
        .ZN(n2077) );
  AOI22_X1 U1395 ( .A1(n2843), .A2(\bank_register[26][3] ), .B1(n2832), .B2(
        \bank_register[14][3] ), .ZN(n2079) );
  OAI21_X1 U1396 ( .B1(n2051), .B2(n2052), .A(n2916), .ZN(n2050) );
  OAI221_X1 U1397 ( .B1(n920), .B2(n2865), .C1(n919), .C2(n2854), .A(n2054), 
        .ZN(n2051) );
  OAI221_X1 U1398 ( .B1(n916), .B2(n2909), .C1(n915), .C2(n2898), .A(n2053), 
        .ZN(n2052) );
  AOI22_X1 U1399 ( .A1(n2843), .A2(\bank_register[26][4] ), .B1(n2832), .B2(
        \bank_register[14][4] ), .ZN(n2054) );
  OAI21_X1 U1400 ( .B1(n2026), .B2(n2027), .A(n2916), .ZN(n2025) );
  OAI221_X1 U1401 ( .B1(n883), .B2(n2865), .C1(n882), .C2(n2854), .A(n2029), 
        .ZN(n2026) );
  OAI221_X1 U1402 ( .B1(n879), .B2(n2909), .C1(n878), .C2(n2898), .A(n2028), 
        .ZN(n2027) );
  AOI22_X1 U1403 ( .A1(n2842), .A2(\bank_register[26][5] ), .B1(n2832), .B2(
        \bank_register[14][5] ), .ZN(n2029) );
  OAI21_X1 U1404 ( .B1(n1951), .B2(n1952), .A(n2916), .ZN(n1950) );
  OAI221_X1 U1405 ( .B1(n772), .B2(n2866), .C1(n771), .C2(n2855), .A(n1954), 
        .ZN(n1951) );
  OAI221_X1 U1406 ( .B1(n768), .B2(n2909), .C1(n767), .C2(n2899), .A(n1953), 
        .ZN(n1952) );
  AOI22_X1 U1407 ( .A1(n2842), .A2(\bank_register[26][8] ), .B1(n2833), .B2(
        \bank_register[14][8] ), .ZN(n1954) );
  OAI21_X1 U1408 ( .B1(n1908), .B2(n1909), .A(n2916), .ZN(n1907) );
  OAI221_X1 U1409 ( .B1(n735), .B2(n2866), .C1(n734), .C2(n2855), .A(n1918), 
        .ZN(n1908) );
  OAI221_X1 U1410 ( .B1(n731), .B2(n2910), .C1(n730), .C2(n2899), .A(n1913), 
        .ZN(n1909) );
  AOI22_X1 U1411 ( .A1(n2844), .A2(\bank_register[26][9] ), .B1(n2833), .B2(
        \bank_register[14][9] ), .ZN(n1918) );
  OAI21_X1 U1412 ( .B1(n2439), .B2(n2440), .A(n2915), .ZN(n2438) );
  OAI221_X1 U1413 ( .B1(n1401), .B2(n2867), .C1(n1400), .C2(n2856), .A(n2442), 
        .ZN(n2439) );
  OAI221_X1 U1414 ( .B1(n1397), .B2(n2911), .C1(n1396), .C2(n2900), .A(n2441), 
        .ZN(n2440) );
  AOI22_X1 U1415 ( .A1(n2845), .A2(\bank_register[26][21] ), .B1(n2834), .B2(
        \bank_register[14][21] ), .ZN(n2442) );
  OAI21_X1 U1416 ( .B1(n2414), .B2(n2415), .A(n2915), .ZN(n2413) );
  OAI221_X1 U1417 ( .B1(n1364), .B2(n2867), .C1(n1363), .C2(n2856), .A(n2417), 
        .ZN(n2414) );
  OAI221_X1 U1418 ( .B1(n1360), .B2(n2911), .C1(n1359), .C2(n2900), .A(n2416), 
        .ZN(n2415) );
  AOI22_X1 U1419 ( .A1(n2845), .A2(\bank_register[26][22] ), .B1(n2834), .B2(
        \bank_register[14][22] ), .ZN(n2417) );
  OAI21_X1 U1420 ( .B1(n2389), .B2(n2390), .A(n2915), .ZN(n2388) );
  OAI221_X1 U1421 ( .B1(n1327), .B2(n2867), .C1(n1326), .C2(n2856), .A(n2392), 
        .ZN(n2389) );
  OAI221_X1 U1422 ( .B1(n1323), .B2(n2911), .C1(n1322), .C2(n2900), .A(n2391), 
        .ZN(n2390) );
  AOI22_X1 U1423 ( .A1(n2845), .A2(\bank_register[26][23] ), .B1(n2834), .B2(
        \bank_register[14][23] ), .ZN(n2392) );
  OAI21_X1 U1424 ( .B1(n2362), .B2(n2363), .A(n2915), .ZN(n2360) );
  OAI221_X1 U1425 ( .B1(n1290), .B2(n2867), .C1(n1289), .C2(n2856), .A(n2366), 
        .ZN(n2362) );
  OAI221_X1 U1426 ( .B1(n1286), .B2(n2911), .C1(n1285), .C2(n2900), .A(n2364), 
        .ZN(n2363) );
  AOI22_X1 U1427 ( .A1(n2845), .A2(\bank_register[26][24] ), .B1(n2834), .B2(
        \bank_register[14][24] ), .ZN(n2366) );
  OAI21_X1 U1428 ( .B1(n2328), .B2(n2330), .A(n2915), .ZN(n2327) );
  OAI221_X1 U1429 ( .B1(n1253), .B2(n2867), .C1(n1252), .C2(n2856), .A(n2332), 
        .ZN(n2328) );
  OAI221_X1 U1430 ( .B1(n1249), .B2(n2910), .C1(n1248), .C2(n2900), .A(n2331), 
        .ZN(n2330) );
  AOI22_X1 U1431 ( .A1(n2845), .A2(\bank_register[26][25] ), .B1(n2834), .B2(
        \bank_register[14][25] ), .ZN(n2332) );
  OAI21_X1 U1432 ( .B1(n2295), .B2(n2296), .A(n2915), .ZN(n2294) );
  OAI221_X1 U1433 ( .B1(n1216), .B2(n2866), .C1(n1215), .C2(n2856), .A(n2299), 
        .ZN(n2295) );
  OAI221_X1 U1434 ( .B1(n1212), .B2(n2910), .C1(n1211), .C2(n2900), .A(n2298), 
        .ZN(n2296) );
  AOI22_X1 U1435 ( .A1(n2844), .A2(\bank_register[26][26] ), .B1(n2834), .B2(
        \bank_register[14][26] ), .ZN(n2299) );
  OAI21_X1 U1436 ( .B1(n2262), .B2(n2263), .A(n2915), .ZN(n2260) );
  OAI221_X1 U1437 ( .B1(n1179), .B2(n2866), .C1(n1178), .C2(n2855), .A(n2266), 
        .ZN(n2262) );
  OAI221_X1 U1438 ( .B1(n1175), .B2(n2910), .C1(n1174), .C2(n2899), .A(n2264), 
        .ZN(n2263) );
  AOI22_X1 U1439 ( .A1(n2844), .A2(\bank_register[26][27] ), .B1(n2833), .B2(
        \bank_register[14][27] ), .ZN(n2266) );
  OAI21_X1 U1440 ( .B1(n2226), .B2(n2228), .A(n2915), .ZN(n2225) );
  OAI221_X1 U1441 ( .B1(n1142), .B2(n2866), .C1(n1141), .C2(n2855), .A(n2231), 
        .ZN(n2226) );
  OAI221_X1 U1442 ( .B1(n1138), .B2(n2910), .C1(n1137), .C2(n2899), .A(n2229), 
        .ZN(n2228) );
  AOI22_X1 U1443 ( .A1(n2844), .A2(\bank_register[26][28] ), .B1(n2833), .B2(
        \bank_register[14][28] ), .ZN(n2231) );
  OAI21_X1 U1444 ( .B1(n2189), .B2(n2190), .A(n2915), .ZN(n2187) );
  OAI221_X1 U1445 ( .B1(n1105), .B2(n2866), .C1(n1104), .C2(n2855), .A(n2193), 
        .ZN(n2189) );
  OAI221_X1 U1446 ( .B1(n1101), .B2(n2909), .C1(n1100), .C2(n2899), .A(n2192), 
        .ZN(n2190) );
  AOI22_X1 U1447 ( .A1(n2844), .A2(\bank_register[26][29] ), .B1(n2833), .B2(
        \bank_register[14][29] ), .ZN(n2193) );
  OAI21_X1 U1448 ( .B1(n2126), .B2(n2127), .A(n2915), .ZN(n2125) );
  OAI221_X1 U1449 ( .B1(n1031), .B2(n2865), .C1(n1030), .C2(n2854), .A(n2129), 
        .ZN(n2126) );
  OAI221_X1 U1450 ( .B1(n1027), .B2(n2909), .C1(n1026), .C2(n2898), .A(n2128), 
        .ZN(n2127) );
  AOI22_X1 U1451 ( .A1(n2843), .A2(\bank_register[26][30] ), .B1(n2832), .B2(
        \bank_register[14][30] ), .ZN(n2129) );
  OAI21_X1 U1452 ( .B1(n2101), .B2(n2102), .A(n2916), .ZN(n2100) );
  OAI221_X1 U1453 ( .B1(n994), .B2(n2866), .C1(n993), .C2(n2855), .A(n2104), 
        .ZN(n2101) );
  OAI221_X1 U1454 ( .B1(n990), .B2(n2910), .C1(n989), .C2(n2899), .A(n2103), 
        .ZN(n2102) );
  AOI22_X1 U1455 ( .A1(n2843), .A2(\bank_register[26][31] ), .B1(n2833), .B2(
        \bank_register[14][31] ), .ZN(n2104) );
  OAI21_X1 U1456 ( .B1(n2489), .B2(n2490), .A(n2914), .ZN(n2488) );
  OAI221_X1 U1457 ( .B1(n1475), .B2(n2867), .C1(n1474), .C2(n2857), .A(n2492), 
        .ZN(n2489) );
  OAI221_X1 U1458 ( .B1(n1471), .B2(n2911), .C1(n1470), .C2(n2901), .A(n2491), 
        .ZN(n2490) );
  AOI22_X1 U1459 ( .A1(n2846), .A2(\bank_register[26][1] ), .B1(n2835), .B2(
        \bank_register[14][1] ), .ZN(n2492) );
  OAI21_X1 U1460 ( .B1(n2664), .B2(n2665), .A(n2914), .ZN(n2663) );
  OAI221_X1 U1461 ( .B1(n1734), .B2(n2869), .C1(n1733), .C2(n2858), .A(n2667), 
        .ZN(n2664) );
  OAI221_X1 U1462 ( .B1(n1730), .B2(n2912), .C1(n1729), .C2(n2902), .A(n2666), 
        .ZN(n2665) );
  AOI22_X1 U1463 ( .A1(n2847), .A2(\bank_register[26][13] ), .B1(n2836), .B2(
        \bank_register[14][13] ), .ZN(n2667) );
  OAI21_X1 U1464 ( .B1(n2639), .B2(n2640), .A(n2914), .ZN(n2638) );
  OAI221_X1 U1465 ( .B1(n1697), .B2(n2868), .C1(n1696), .C2(n2858), .A(n2642), 
        .ZN(n2639) );
  OAI221_X1 U1466 ( .B1(n1693), .B2(n2912), .C1(n1692), .C2(n2902), .A(n2641), 
        .ZN(n2640) );
  AOI22_X1 U1467 ( .A1(n2847), .A2(\bank_register[26][14] ), .B1(n2836), .B2(
        \bank_register[14][14] ), .ZN(n2642) );
  OAI21_X1 U1468 ( .B1(n2614), .B2(n2615), .A(n2914), .ZN(n2613) );
  OAI221_X1 U1469 ( .B1(n1660), .B2(n2868), .C1(n1659), .C2(n2858), .A(n2617), 
        .ZN(n2614) );
  OAI221_X1 U1470 ( .B1(n1656), .B2(n2912), .C1(n1655), .C2(n2902), .A(n2616), 
        .ZN(n2615) );
  AOI22_X1 U1471 ( .A1(n2846), .A2(\bank_register[26][15] ), .B1(n2836), .B2(
        \bank_register[14][15] ), .ZN(n2617) );
  OAI21_X1 U1472 ( .B1(n2589), .B2(n2590), .A(n2914), .ZN(n2588) );
  OAI221_X1 U1473 ( .B1(n1623), .B2(n2868), .C1(n1622), .C2(n2857), .A(n2592), 
        .ZN(n2589) );
  OAI221_X1 U1474 ( .B1(n1619), .B2(n2912), .C1(n1618), .C2(n2901), .A(n2591), 
        .ZN(n2590) );
  AOI22_X1 U1475 ( .A1(n2846), .A2(\bank_register[26][16] ), .B1(n2835), .B2(
        \bank_register[14][16] ), .ZN(n2592) );
  OAI21_X1 U1476 ( .B1(n2564), .B2(n2565), .A(n2914), .ZN(n2563) );
  OAI221_X1 U1477 ( .B1(n1586), .B2(n2868), .C1(n1585), .C2(n2857), .A(n2567), 
        .ZN(n2564) );
  OAI221_X1 U1478 ( .B1(n1582), .B2(n2912), .C1(n1581), .C2(n2901), .A(n2566), 
        .ZN(n2565) );
  AOI22_X1 U1479 ( .A1(n2846), .A2(\bank_register[26][17] ), .B1(n2835), .B2(
        \bank_register[14][17] ), .ZN(n2567) );
  OAI21_X1 U1480 ( .B1(n2539), .B2(n2540), .A(n2914), .ZN(n2538) );
  OAI221_X1 U1481 ( .B1(n1549), .B2(n2868), .C1(n1548), .C2(n2857), .A(n2542), 
        .ZN(n2539) );
  OAI221_X1 U1482 ( .B1(n1545), .B2(n2912), .C1(n1544), .C2(n2901), .A(n2541), 
        .ZN(n2540) );
  AOI22_X1 U1483 ( .A1(n2846), .A2(\bank_register[26][18] ), .B1(n2835), .B2(
        \bank_register[14][18] ), .ZN(n2542) );
  OAI21_X1 U1484 ( .B1(n2514), .B2(n2515), .A(n2914), .ZN(n2513) );
  OAI221_X1 U1485 ( .B1(n1512), .B2(n2868), .C1(n1511), .C2(n2857), .A(n2517), 
        .ZN(n2514) );
  OAI221_X1 U1486 ( .B1(n1508), .B2(n2912), .C1(n1507), .C2(n2901), .A(n2516), 
        .ZN(n2515) );
  AOI22_X1 U1487 ( .A1(n2846), .A2(\bank_register[26][19] ), .B1(n2835), .B2(
        \bank_register[14][19] ), .ZN(n2517) );
  OAI21_X1 U1488 ( .B1(n2464), .B2(n2465), .A(n2915), .ZN(n2463) );
  OAI221_X1 U1489 ( .B1(n1438), .B2(n2867), .C1(n1437), .C2(n2857), .A(n2467), 
        .ZN(n2464) );
  OAI221_X1 U1490 ( .B1(n1434), .B2(n2911), .C1(n1433), .C2(n2901), .A(n2466), 
        .ZN(n2465) );
  AOI22_X1 U1491 ( .A1(n2845), .A2(\bank_register[26][20] ), .B1(n2835), .B2(
        \bank_register[14][20] ), .ZN(n2467) );
  INV_X1 U1492 ( .A(read_address_2[3]), .ZN(n1888) );
  INV_X1 U1493 ( .A(read_address_1[2]), .ZN(n2787) );
  OAI21_X1 U1494 ( .B1(n2775), .B2(n2776), .A(n2820), .ZN(n2761) );
  OAI221_X1 U1495 ( .B1(n2790), .B2(n2808), .C1(n2791), .C2(n2805), .A(n2792), 
        .ZN(n2775) );
  OAI221_X1 U1496 ( .B1(n2777), .B2(n2817), .C1(n2778), .C2(n2814), .A(n2779), 
        .ZN(n2776) );
  INV_X1 U1497 ( .A(\bank_register[12][0] ), .ZN(n2791) );
  OAI21_X1 U1498 ( .B1(n2497), .B2(n2498), .A(n2820), .ZN(n2486) );
  OAI221_X1 U1499 ( .B1(n2507), .B2(n2808), .C1(n2508), .C2(n2805), .A(n2509), 
        .ZN(n2497) );
  OAI221_X1 U1500 ( .B1(n2499), .B2(n2817), .C1(n2500), .C2(n2814), .A(n2501), 
        .ZN(n2498) );
  INV_X1 U1501 ( .A(\bank_register[12][1] ), .ZN(n2508) );
  OAI21_X1 U1502 ( .B1(n2163), .B2(n2165), .A(n2821), .ZN(n2148) );
  OAI221_X1 U1503 ( .B1(n2178), .B2(n2809), .C1(n2180), .C2(n2806), .A(n2181), 
        .ZN(n2163) );
  OAI221_X1 U1504 ( .B1(n2166), .B2(n2818), .C1(n2168), .C2(n2815), .A(n2169), 
        .ZN(n2165) );
  INV_X1 U1505 ( .A(\bank_register[12][2] ), .ZN(n2180) );
  OAI21_X1 U1506 ( .B1(n2747), .B2(n2748), .A(n2820), .ZN(n2736) );
  OAI221_X1 U1507 ( .B1(n2757), .B2(n2808), .C1(n2758), .C2(n2805), .A(n2759), 
        .ZN(n2747) );
  OAI221_X1 U1508 ( .B1(n2749), .B2(n2817), .C1(n2750), .C2(n2814), .A(n2751), 
        .ZN(n2748) );
  INV_X1 U1509 ( .A(\bank_register[12][10] ), .ZN(n2758) );
  OAI21_X1 U1510 ( .B1(n2722), .B2(n2723), .A(n2820), .ZN(n2711) );
  OAI221_X1 U1511 ( .B1(n2732), .B2(n2808), .C1(n2733), .C2(n2805), .A(n2734), 
        .ZN(n2722) );
  OAI221_X1 U1512 ( .B1(n2724), .B2(n2817), .C1(n2725), .C2(n2814), .A(n2726), 
        .ZN(n2723) );
  INV_X1 U1513 ( .A(\bank_register[12][11] ), .ZN(n2733) );
  OAI21_X1 U1514 ( .B1(n2697), .B2(n2698), .A(n2820), .ZN(n2686) );
  OAI221_X1 U1515 ( .B1(n2707), .B2(n2808), .C1(n2708), .C2(n2805), .A(n2709), 
        .ZN(n2697) );
  OAI221_X1 U1516 ( .B1(n2699), .B2(n2817), .C1(n2700), .C2(n2814), .A(n2701), 
        .ZN(n2698) );
  INV_X1 U1517 ( .A(\bank_register[12][12] ), .ZN(n2708) );
  OAI21_X1 U1518 ( .B1(n2672), .B2(n2673), .A(n2820), .ZN(n2661) );
  OAI221_X1 U1519 ( .B1(n2682), .B2(n2808), .C1(n2683), .C2(n2805), .A(n2684), 
        .ZN(n2672) );
  OAI221_X1 U1520 ( .B1(n2674), .B2(n2817), .C1(n2675), .C2(n2814), .A(n2676), 
        .ZN(n2673) );
  INV_X1 U1521 ( .A(\bank_register[12][13] ), .ZN(n2683) );
  OAI21_X1 U1522 ( .B1(n2647), .B2(n2648), .A(n2820), .ZN(n2636) );
  OAI221_X1 U1523 ( .B1(n2657), .B2(n2808), .C1(n2658), .C2(n2805), .A(n2659), 
        .ZN(n2647) );
  OAI221_X1 U1524 ( .B1(n2649), .B2(n2817), .C1(n2650), .C2(n2814), .A(n2651), 
        .ZN(n2648) );
  INV_X1 U1525 ( .A(\bank_register[12][14] ), .ZN(n2658) );
  OAI21_X1 U1526 ( .B1(n2622), .B2(n2623), .A(n2820), .ZN(n2611) );
  OAI221_X1 U1527 ( .B1(n2632), .B2(n2808), .C1(n2633), .C2(n2805), .A(n2634), 
        .ZN(n2622) );
  OAI221_X1 U1528 ( .B1(n2624), .B2(n2817), .C1(n2625), .C2(n2814), .A(n2626), 
        .ZN(n2623) );
  INV_X1 U1529 ( .A(\bank_register[12][15] ), .ZN(n2633) );
  OAI21_X1 U1530 ( .B1(n2597), .B2(n2598), .A(n2820), .ZN(n2586) );
  OAI221_X1 U1531 ( .B1(n2607), .B2(n2808), .C1(n2608), .C2(n2805), .A(n2609), 
        .ZN(n2597) );
  OAI221_X1 U1532 ( .B1(n2599), .B2(n2817), .C1(n2600), .C2(n2814), .A(n2601), 
        .ZN(n2598) );
  INV_X1 U1533 ( .A(\bank_register[12][16] ), .ZN(n2608) );
  OAI21_X1 U1534 ( .B1(n2572), .B2(n2573), .A(n2820), .ZN(n2561) );
  OAI221_X1 U1535 ( .B1(n2582), .B2(n2808), .C1(n2583), .C2(n2805), .A(n2584), 
        .ZN(n2572) );
  OAI221_X1 U1536 ( .B1(n2574), .B2(n2817), .C1(n2575), .C2(n2814), .A(n2576), 
        .ZN(n2573) );
  INV_X1 U1537 ( .A(\bank_register[12][17] ), .ZN(n2583) );
  OAI21_X1 U1538 ( .B1(n2547), .B2(n2548), .A(n2820), .ZN(n2536) );
  OAI221_X1 U1539 ( .B1(n2557), .B2(n2808), .C1(n2558), .C2(n2805), .A(n2559), 
        .ZN(n2547) );
  OAI221_X1 U1540 ( .B1(n2549), .B2(n2817), .C1(n2550), .C2(n2814), .A(n2551), 
        .ZN(n2548) );
  INV_X1 U1541 ( .A(\bank_register[12][18] ), .ZN(n2558) );
  OAI21_X1 U1542 ( .B1(n2522), .B2(n2523), .A(n2820), .ZN(n2511) );
  OAI221_X1 U1543 ( .B1(n2532), .B2(n2808), .C1(n2533), .C2(n2805), .A(n2534), 
        .ZN(n2522) );
  OAI221_X1 U1544 ( .B1(n2524), .B2(n2817), .C1(n2525), .C2(n2814), .A(n2526), 
        .ZN(n2523) );
  INV_X1 U1545 ( .A(\bank_register[12][19] ), .ZN(n2533) );
  OAI21_X1 U1546 ( .B1(n2472), .B2(n2473), .A(n2821), .ZN(n2461) );
  OAI221_X1 U1547 ( .B1(n2482), .B2(n2809), .C1(n2483), .C2(n2806), .A(n2484), 
        .ZN(n2472) );
  OAI221_X1 U1548 ( .B1(n2474), .B2(n2818), .C1(n2475), .C2(n2815), .A(n2476), 
        .ZN(n2473) );
  INV_X1 U1549 ( .A(\bank_register[12][20] ), .ZN(n2483) );
  OAI21_X1 U1550 ( .B1(n2447), .B2(n2448), .A(n2821), .ZN(n2436) );
  OAI221_X1 U1551 ( .B1(n2457), .B2(n2809), .C1(n2458), .C2(n2806), .A(n2459), 
        .ZN(n2447) );
  OAI221_X1 U1552 ( .B1(n2449), .B2(n2818), .C1(n2450), .C2(n2815), .A(n2451), 
        .ZN(n2448) );
  INV_X1 U1553 ( .A(\bank_register[12][21] ), .ZN(n2458) );
  OAI21_X1 U1554 ( .B1(n2422), .B2(n2423), .A(n2821), .ZN(n2411) );
  OAI221_X1 U1555 ( .B1(n2432), .B2(n2809), .C1(n2433), .C2(n2806), .A(n2434), 
        .ZN(n2422) );
  OAI221_X1 U1556 ( .B1(n2424), .B2(n2818), .C1(n2425), .C2(n2815), .A(n2426), 
        .ZN(n2423) );
  INV_X1 U1557 ( .A(\bank_register[12][22] ), .ZN(n2433) );
  OAI21_X1 U1558 ( .B1(n2397), .B2(n2398), .A(n2821), .ZN(n2386) );
  OAI221_X1 U1559 ( .B1(n2407), .B2(n2809), .C1(n2408), .C2(n2806), .A(n2409), 
        .ZN(n2397) );
  OAI221_X1 U1560 ( .B1(n2399), .B2(n2818), .C1(n2400), .C2(n2815), .A(n2401), 
        .ZN(n2398) );
  INV_X1 U1561 ( .A(\bank_register[12][23] ), .ZN(n2408) );
  OAI21_X1 U1562 ( .B1(n2372), .B2(n2373), .A(n2821), .ZN(n2358) );
  OAI221_X1 U1563 ( .B1(n2382), .B2(n2809), .C1(n2383), .C2(n2806), .A(n2384), 
        .ZN(n2372) );
  OAI221_X1 U1564 ( .B1(n2374), .B2(n2818), .C1(n2375), .C2(n2815), .A(n2376), 
        .ZN(n2373) );
  INV_X1 U1565 ( .A(\bank_register[12][24] ), .ZN(n2383) );
  OAI21_X1 U1566 ( .B1(n2339), .B2(n2340), .A(n2821), .ZN(n2324) );
  OAI221_X1 U1567 ( .B1(n2352), .B2(n2809), .C1(n2354), .C2(n2806), .A(n2355), 
        .ZN(n2339) );
  OAI221_X1 U1568 ( .B1(n2342), .B2(n2818), .C1(n2343), .C2(n2815), .A(n2344), 
        .ZN(n2340) );
  INV_X1 U1569 ( .A(\bank_register[12][25] ), .ZN(n2354) );
  OAI21_X1 U1570 ( .B1(n2306), .B2(n2307), .A(n2821), .ZN(n2291) );
  OAI221_X1 U1571 ( .B1(n2319), .B2(n2809), .C1(n2320), .C2(n2806), .A(n2322), 
        .ZN(n2306) );
  OAI221_X1 U1572 ( .B1(n2308), .B2(n2818), .C1(n2310), .C2(n2815), .A(n2311), 
        .ZN(n2307) );
  INV_X1 U1573 ( .A(\bank_register[12][26] ), .ZN(n2320) );
  OAI21_X1 U1574 ( .B1(n2272), .B2(n2274), .A(n2821), .ZN(n2258) );
  OAI221_X1 U1575 ( .B1(n2286), .B2(n2809), .C1(n2287), .C2(n2806), .A(n2288), 
        .ZN(n2272) );
  OAI221_X1 U1576 ( .B1(n2275), .B2(n2818), .C1(n2276), .C2(n2815), .A(n2278), 
        .ZN(n2274) );
  INV_X1 U1577 ( .A(\bank_register[12][27] ), .ZN(n2287) );
  OAI21_X1 U1578 ( .B1(n2238), .B2(n2240), .A(n2821), .ZN(n2222) );
  OAI221_X1 U1579 ( .B1(n2252), .B2(n2809), .C1(n2254), .C2(n2806), .A(n2255), 
        .ZN(n2238) );
  OAI221_X1 U1580 ( .B1(n2241), .B2(n2818), .C1(n2243), .C2(n2815), .A(n2244), 
        .ZN(n2240) );
  INV_X1 U1581 ( .A(\bank_register[12][28] ), .ZN(n2254) );
  OAI21_X1 U1582 ( .B1(n2201), .B2(n2202), .A(n2821), .ZN(n2184) );
  OAI221_X1 U1583 ( .B1(n2216), .B2(n2809), .C1(n2217), .C2(n2806), .A(n2219), 
        .ZN(n2201) );
  OAI221_X1 U1584 ( .B1(n2204), .B2(n2818), .C1(n2205), .C2(n2815), .A(n2207), 
        .ZN(n2202) );
  INV_X1 U1585 ( .A(\bank_register[12][29] ), .ZN(n2217) );
  OAI21_X1 U1586 ( .B1(n2134), .B2(n2135), .A(n2821), .ZN(n2123) );
  OAI221_X1 U1587 ( .B1(n2144), .B2(n2809), .C1(n2145), .C2(n2806), .A(n2146), 
        .ZN(n2134) );
  OAI221_X1 U1588 ( .B1(n2136), .B2(n2818), .C1(n2137), .C2(n2815), .A(n2138), 
        .ZN(n2135) );
  INV_X1 U1589 ( .A(\bank_register[12][30] ), .ZN(n2145) );
  OAI21_X1 U1590 ( .B1(n2109), .B2(n2110), .A(n2822), .ZN(n2098) );
  OAI221_X1 U1591 ( .B1(n2119), .B2(n2810), .C1(n2120), .C2(n2807), .A(n2121), 
        .ZN(n2109) );
  OAI221_X1 U1592 ( .B1(n2111), .B2(n2819), .C1(n2112), .C2(n2816), .A(n2113), 
        .ZN(n2110) );
  INV_X1 U1593 ( .A(\bank_register[12][31] ), .ZN(n2120) );
  NAND2_X1 U1594 ( .A1(n1899), .A2(read_address_2[2]), .ZN(n1856) );
  NAND2_X1 U1595 ( .A1(n1898), .A2(read_address_2[2]), .ZN(n1857) );
  NAND2_X1 U1596 ( .A1(n1901), .A2(read_address_2[2]), .ZN(n1854) );
  INV_X1 U1597 ( .A(read_address_2[4]), .ZN(n1895) );
  AOI22_X1 U1598 ( .A1(\bank_register[4][1] ), .A2(n3009), .B1(n3238), .B2(
        n1447), .ZN(n1443) );
  NAND2_X1 U1599 ( .A1(n1448), .A2(n1449), .ZN(n1447) );
  AOI221_X1 U1600 ( .B1(\bank_register[21][1] ), .B2(n2957), .C1(
        \bank_register[29][1] ), .C2(n2946), .A(n1453), .ZN(n1448) );
  AOI221_X1 U1601 ( .B1(\bank_register[25][1] ), .B2(n3001), .C1(
        \bank_register[13][1] ), .C2(n2990), .A(n1450), .ZN(n1449) );
  AOI22_X1 U1602 ( .A1(\bank_register[4][2] ), .A2(n3010), .B1(n3238), .B2(
        n1040), .ZN(n1036) );
  NAND2_X1 U1603 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
  AOI221_X1 U1604 ( .B1(\bank_register[21][2] ), .B2(n2956), .C1(
        \bank_register[29][2] ), .C2(n2945), .A(n1046), .ZN(n1041) );
  AOI221_X1 U1605 ( .B1(\bank_register[25][2] ), .B2(n3000), .C1(
        \bank_register[13][2] ), .C2(n2989), .A(n1043), .ZN(n1042) );
  AOI22_X1 U1606 ( .A1(\bank_register[4][3] ), .A2(n3011), .B1(n3238), .B2(
        n929), .ZN(n925) );
  NAND2_X1 U1607 ( .A1(n930), .A2(n931), .ZN(n929) );
  AOI221_X1 U1608 ( .B1(\bank_register[21][3] ), .B2(n2956), .C1(
        \bank_register[29][3] ), .C2(n2945), .A(n935), .ZN(n930) );
  AOI221_X1 U1609 ( .B1(\bank_register[25][3] ), .B2(n3000), .C1(
        \bank_register[13][3] ), .C2(n2989), .A(n932), .ZN(n931) );
  AOI22_X1 U1610 ( .A1(\bank_register[4][4] ), .A2(n3011), .B1(n3238), .B2(
        n892), .ZN(n888) );
  NAND2_X1 U1611 ( .A1(n893), .A2(n894), .ZN(n892) );
  AOI221_X1 U1612 ( .B1(\bank_register[21][4] ), .B2(n2956), .C1(
        \bank_register[29][4] ), .C2(n2945), .A(n898), .ZN(n893) );
  AOI221_X1 U1613 ( .B1(\bank_register[25][4] ), .B2(n3000), .C1(
        \bank_register[13][4] ), .C2(n2989), .A(n895), .ZN(n894) );
  AOI22_X1 U1614 ( .A1(\bank_register[4][5] ), .A2(n3011), .B1(n3238), .B2(
        n855), .ZN(n851) );
  NAND2_X1 U1615 ( .A1(n856), .A2(n857), .ZN(n855) );
  AOI221_X1 U1616 ( .B1(\bank_register[21][5] ), .B2(n2956), .C1(
        \bank_register[29][5] ), .C2(n2945), .A(n861), .ZN(n856) );
  AOI221_X1 U1617 ( .B1(\bank_register[25][5] ), .B2(n3000), .C1(
        \bank_register[13][5] ), .C2(n2989), .A(n858), .ZN(n857) );
  AOI22_X1 U1618 ( .A1(\bank_register[4][6] ), .A2(n3011), .B1(
        read_address_2[0]), .B2(n818), .ZN(n814) );
  NAND2_X1 U1619 ( .A1(n819), .A2(n820), .ZN(n818) );
  AOI221_X1 U1620 ( .B1(\bank_register[21][6] ), .B2(n2956), .C1(
        \bank_register[29][6] ), .C2(n2945), .A(n824), .ZN(n819) );
  AOI221_X1 U1621 ( .B1(\bank_register[25][6] ), .B2(n3000), .C1(
        \bank_register[13][6] ), .C2(n2989), .A(n821), .ZN(n820) );
  AOI22_X1 U1622 ( .A1(\bank_register[4][7] ), .A2(n3011), .B1(
        read_address_2[0]), .B2(n781), .ZN(n777) );
  NAND2_X1 U1623 ( .A1(n782), .A2(n783), .ZN(n781) );
  AOI221_X1 U1624 ( .B1(\bank_register[21][7] ), .B2(n2956), .C1(
        \bank_register[29][7] ), .C2(n2945), .A(n787), .ZN(n782) );
  AOI221_X1 U1625 ( .B1(\bank_register[25][7] ), .B2(n3000), .C1(
        \bank_register[13][7] ), .C2(n2989), .A(n784), .ZN(n783) );
  AOI22_X1 U1626 ( .A1(\bank_register[4][8] ), .A2(n3011), .B1(
        read_address_2[0]), .B2(n744), .ZN(n740) );
  NAND2_X1 U1627 ( .A1(n745), .A2(n746), .ZN(n744) );
  AOI221_X1 U1628 ( .B1(\bank_register[21][8] ), .B2(n2956), .C1(
        \bank_register[29][8] ), .C2(n2945), .A(n750), .ZN(n745) );
  AOI221_X1 U1629 ( .B1(\bank_register[25][8] ), .B2(n3000), .C1(
        \bank_register[13][8] ), .C2(n2989), .A(n747), .ZN(n746) );
  AOI22_X1 U1630 ( .A1(\bank_register[4][9] ), .A2(n3011), .B1(
        read_address_2[0]), .B2(n699), .ZN(n688) );
  NAND2_X1 U1631 ( .A1(n700), .A2(n701), .ZN(n699) );
  AOI221_X1 U1632 ( .B1(\bank_register[21][9] ), .B2(n2957), .C1(
        \bank_register[29][9] ), .C2(n2946), .A(n711), .ZN(n700) );
  AOI221_X1 U1633 ( .B1(\bank_register[25][9] ), .B2(n3001), .C1(
        \bank_register[13][9] ), .C2(n2990), .A(n704), .ZN(n701) );
  AOI22_X1 U1634 ( .A1(\bank_register[4][17] ), .A2(n3009), .B1(n3238), .B2(
        n1558), .ZN(n1554) );
  NAND2_X1 U1635 ( .A1(n1559), .A2(n1560), .ZN(n1558) );
  AOI221_X1 U1636 ( .B1(\bank_register[21][17] ), .B2(n2957), .C1(
        \bank_register[29][17] ), .C2(n2946), .A(n1564), .ZN(n1559) );
  AOI221_X1 U1637 ( .B1(\bank_register[25][17] ), .B2(n3001), .C1(
        \bank_register[13][17] ), .C2(n2990), .A(n1561), .ZN(n1560) );
  AOI22_X1 U1638 ( .A1(\bank_register[4][18] ), .A2(n3009), .B1(n3238), .B2(
        n1521), .ZN(n1517) );
  NAND2_X1 U1639 ( .A1(n1522), .A2(n1523), .ZN(n1521) );
  AOI221_X1 U1640 ( .B1(\bank_register[21][18] ), .B2(n2957), .C1(
        \bank_register[29][18] ), .C2(n2946), .A(n1527), .ZN(n1522) );
  AOI221_X1 U1641 ( .B1(\bank_register[25][18] ), .B2(n3001), .C1(
        \bank_register[13][18] ), .C2(n2990), .A(n1524), .ZN(n1523) );
  AOI22_X1 U1642 ( .A1(\bank_register[4][19] ), .A2(n3009), .B1(n3238), .B2(
        n1484), .ZN(n1480) );
  NAND2_X1 U1643 ( .A1(n1485), .A2(n1486), .ZN(n1484) );
  AOI221_X1 U1644 ( .B1(\bank_register[21][19] ), .B2(n2957), .C1(
        \bank_register[29][19] ), .C2(n2946), .A(n1490), .ZN(n1485) );
  AOI221_X1 U1645 ( .B1(\bank_register[25][19] ), .B2(n3001), .C1(
        \bank_register[13][19] ), .C2(n2990), .A(n1487), .ZN(n1486) );
  AOI22_X1 U1646 ( .A1(\bank_register[4][20] ), .A2(n3010), .B1(n3238), .B2(
        n1410), .ZN(n1406) );
  NAND2_X1 U1647 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
  AOI221_X1 U1648 ( .B1(\bank_register[21][20] ), .B2(n2957), .C1(
        \bank_register[29][20] ), .C2(n2946), .A(n1416), .ZN(n1411) );
  AOI221_X1 U1649 ( .B1(\bank_register[25][20] ), .B2(n3001), .C1(
        \bank_register[13][20] ), .C2(n2990), .A(n1413), .ZN(n1412) );
  AOI22_X1 U1650 ( .A1(\bank_register[4][21] ), .A2(n3010), .B1(n3238), .B2(
        n1373), .ZN(n1369) );
  NAND2_X1 U1651 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
  AOI221_X1 U1652 ( .B1(\bank_register[21][21] ), .B2(n2957), .C1(
        \bank_register[29][21] ), .C2(n2946), .A(n1379), .ZN(n1374) );
  AOI221_X1 U1653 ( .B1(\bank_register[25][21] ), .B2(n3001), .C1(
        \bank_register[13][21] ), .C2(n2990), .A(n1376), .ZN(n1375) );
  AOI22_X1 U1654 ( .A1(\bank_register[4][22] ), .A2(n3010), .B1(n3238), .B2(
        n1336), .ZN(n1332) );
  NAND2_X1 U1655 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
  AOI221_X1 U1656 ( .B1(\bank_register[21][22] ), .B2(n2957), .C1(
        \bank_register[29][22] ), .C2(n2946), .A(n1342), .ZN(n1337) );
  AOI221_X1 U1657 ( .B1(\bank_register[25][22] ), .B2(n3001), .C1(
        \bank_register[13][22] ), .C2(n2990), .A(n1339), .ZN(n1338) );
  AOI22_X1 U1658 ( .A1(\bank_register[4][23] ), .A2(n3010), .B1(n3238), .B2(
        n1299), .ZN(n1295) );
  NAND2_X1 U1659 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
  AOI221_X1 U1660 ( .B1(\bank_register[21][23] ), .B2(n2957), .C1(
        \bank_register[29][23] ), .C2(n2946), .A(n1305), .ZN(n1300) );
  AOI221_X1 U1661 ( .B1(\bank_register[25][23] ), .B2(n3001), .C1(
        \bank_register[13][23] ), .C2(n2990), .A(n1302), .ZN(n1301) );
  AOI22_X1 U1662 ( .A1(\bank_register[4][24] ), .A2(n3010), .B1(n3238), .B2(
        n1262), .ZN(n1258) );
  NAND2_X1 U1663 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
  AOI221_X1 U1664 ( .B1(\bank_register[21][24] ), .B2(n2957), .C1(
        \bank_register[29][24] ), .C2(n2946), .A(n1268), .ZN(n1263) );
  AOI221_X1 U1665 ( .B1(\bank_register[25][24] ), .B2(n3001), .C1(
        \bank_register[13][24] ), .C2(n2990), .A(n1265), .ZN(n1264) );
  AOI22_X1 U1666 ( .A1(\bank_register[4][25] ), .A2(n3010), .B1(n3238), .B2(
        n1225), .ZN(n1221) );
  NAND2_X1 U1667 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
  AOI221_X1 U1668 ( .B1(\bank_register[21][25] ), .B2(n2957), .C1(
        \bank_register[29][25] ), .C2(n2946), .A(n1231), .ZN(n1226) );
  AOI221_X1 U1669 ( .B1(\bank_register[25][25] ), .B2(n3001), .C1(
        \bank_register[13][25] ), .C2(n2990), .A(n1228), .ZN(n1227) );
  AOI22_X1 U1670 ( .A1(\bank_register[4][26] ), .A2(n3010), .B1(n3238), .B2(
        n1188), .ZN(n1184) );
  NAND2_X1 U1671 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
  AOI221_X1 U1672 ( .B1(\bank_register[21][26] ), .B2(n2957), .C1(
        \bank_register[29][26] ), .C2(n2946), .A(n1194), .ZN(n1189) );
  AOI221_X1 U1673 ( .B1(\bank_register[25][26] ), .B2(n3001), .C1(
        \bank_register[13][26] ), .C2(n2990), .A(n1191), .ZN(n1190) );
  AOI22_X1 U1674 ( .A1(\bank_register[4][27] ), .A2(n3010), .B1(n3238), .B2(
        n1151), .ZN(n1147) );
  NAND2_X1 U1675 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
  AOI221_X1 U1676 ( .B1(\bank_register[21][27] ), .B2(n2956), .C1(
        \bank_register[29][27] ), .C2(n2945), .A(n1157), .ZN(n1152) );
  AOI221_X1 U1677 ( .B1(\bank_register[25][27] ), .B2(n3000), .C1(
        \bank_register[13][27] ), .C2(n2989), .A(n1154), .ZN(n1153) );
  AOI22_X1 U1678 ( .A1(\bank_register[4][28] ), .A2(n3010), .B1(n3238), .B2(
        n1114), .ZN(n1110) );
  NAND2_X1 U1679 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
  AOI221_X1 U1680 ( .B1(\bank_register[21][28] ), .B2(n2956), .C1(
        \bank_register[29][28] ), .C2(n2945), .A(n1120), .ZN(n1115) );
  AOI221_X1 U1681 ( .B1(\bank_register[25][28] ), .B2(n3000), .C1(
        \bank_register[13][28] ), .C2(n2989), .A(n1117), .ZN(n1116) );
  AOI22_X1 U1682 ( .A1(\bank_register[4][29] ), .A2(n3010), .B1(n3238), .B2(
        n1077), .ZN(n1073) );
  NAND2_X1 U1683 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
  AOI221_X1 U1684 ( .B1(\bank_register[21][29] ), .B2(n2956), .C1(
        \bank_register[29][29] ), .C2(n2945), .A(n1083), .ZN(n1078) );
  AOI221_X1 U1685 ( .B1(\bank_register[25][29] ), .B2(n3000), .C1(
        \bank_register[13][29] ), .C2(n2989), .A(n1080), .ZN(n1079) );
  AOI22_X1 U1686 ( .A1(\bank_register[4][30] ), .A2(n3010), .B1(n3238), .B2(
        n1003), .ZN(n999) );
  NAND2_X1 U1687 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
  AOI221_X1 U1688 ( .B1(\bank_register[21][30] ), .B2(n2956), .C1(
        \bank_register[29][30] ), .C2(n2945), .A(n1009), .ZN(n1004) );
  AOI221_X1 U1689 ( .B1(\bank_register[25][30] ), .B2(n3000), .C1(
        \bank_register[13][30] ), .C2(n2989), .A(n1006), .ZN(n1005) );
  AOI22_X1 U1690 ( .A1(\bank_register[4][31] ), .A2(n3011), .B1(
        read_address_2[0]), .B2(n966), .ZN(n962) );
  NAND2_X1 U1691 ( .A1(n967), .A2(n968), .ZN(n966) );
  AOI221_X1 U1692 ( .B1(\bank_register[21][31] ), .B2(n2956), .C1(
        \bank_register[29][31] ), .C2(n2945), .A(n972), .ZN(n967) );
  AOI221_X1 U1693 ( .B1(\bank_register[25][31] ), .B2(n3000), .C1(
        \bank_register[13][31] ), .C2(n2989), .A(n969), .ZN(n968) );
  INV_X1 U1694 ( .A(read_address_2[1]), .ZN(n1879) );
  INV_X1 U1695 ( .A(n1897), .ZN(n1891) );
  AOI22_X1 U1696 ( .A1(n2952), .A2(\bank_register[30][0] ), .B1(n2963), .B2(
        \bank_register[22][0] ), .ZN(n1897) );
  INV_X1 U1697 ( .A(n1874), .ZN(n1870) );
  AOI22_X1 U1698 ( .A1(n2952), .A2(\bank_register[31][0] ), .B1(n2963), .B2(
        \bank_register[23][0] ), .ZN(n1874) );
  INV_X1 U1699 ( .A(n796), .ZN(n792) );
  AOI22_X1 U1700 ( .A1(n2952), .A2(\bank_register[31][7] ), .B1(n2963), .B2(
        \bank_register[23][7] ), .ZN(n796) );
  INV_X1 U1701 ( .A(n769), .ZN(n765) );
  AOI22_X1 U1702 ( .A1(n2952), .A2(\bank_register[30][8] ), .B1(n2963), .B2(
        \bank_register[22][8] ), .ZN(n769) );
  INV_X1 U1703 ( .A(n759), .ZN(n755) );
  AOI22_X1 U1704 ( .A1(n2952), .A2(\bank_register[31][8] ), .B1(n2963), .B2(
        \bank_register[23][8] ), .ZN(n759) );
  INV_X1 U1705 ( .A(n732), .ZN(n728) );
  AOI22_X1 U1706 ( .A1(n2952), .A2(\bank_register[30][9] ), .B1(n2963), .B2(
        \bank_register[22][9] ), .ZN(n732) );
  INV_X1 U1707 ( .A(n722), .ZN(n718) );
  AOI22_X1 U1708 ( .A1(n2952), .A2(\bank_register[31][9] ), .B1(n2963), .B2(
        \bank_register[23][9] ), .ZN(n722) );
  INV_X1 U1709 ( .A(n1832), .ZN(n1828) );
  AOI22_X1 U1710 ( .A1(n2952), .A2(\bank_register[31][10] ), .B1(n2963), .B2(
        \bank_register[23][10] ), .ZN(n1832) );
  INV_X1 U1711 ( .A(n1900), .ZN(n1890) );
  AOI22_X1 U1712 ( .A1(n2996), .A2(\bank_register[14][0] ), .B1(n3007), .B2(
        \bank_register[26][0] ), .ZN(n1900) );
  INV_X1 U1713 ( .A(n1875), .ZN(n1869) );
  AOI22_X1 U1714 ( .A1(n2996), .A2(\bank_register[15][0] ), .B1(n3007), .B2(
        \bank_register[27][0] ), .ZN(n1875) );
  INV_X1 U1715 ( .A(n797), .ZN(n791) );
  AOI22_X1 U1716 ( .A1(n2996), .A2(\bank_register[15][7] ), .B1(n3007), .B2(
        \bank_register[27][7] ), .ZN(n797) );
  INV_X1 U1717 ( .A(n770), .ZN(n764) );
  AOI22_X1 U1718 ( .A1(n2996), .A2(\bank_register[14][8] ), .B1(n3007), .B2(
        \bank_register[26][8] ), .ZN(n770) );
  INV_X1 U1719 ( .A(n760), .ZN(n754) );
  AOI22_X1 U1720 ( .A1(n2996), .A2(\bank_register[15][8] ), .B1(n3007), .B2(
        \bank_register[27][8] ), .ZN(n760) );
  INV_X1 U1721 ( .A(n733), .ZN(n727) );
  AOI22_X1 U1722 ( .A1(n2996), .A2(\bank_register[14][9] ), .B1(n3007), .B2(
        \bank_register[26][9] ), .ZN(n733) );
  INV_X1 U1723 ( .A(n723), .ZN(n717) );
  AOI22_X1 U1724 ( .A1(n2996), .A2(\bank_register[15][9] ), .B1(n3007), .B2(
        \bank_register[27][9] ), .ZN(n723) );
  INV_X1 U1725 ( .A(n1833), .ZN(n1827) );
  AOI22_X1 U1726 ( .A1(n2996), .A2(\bank_register[15][10] ), .B1(n3007), .B2(
        \bank_register[27][10] ), .ZN(n1833) );
  AND2_X1 U1727 ( .A1(read_address_1[1]), .A2(n2772), .ZN(n2766) );
  AND2_X1 U1728 ( .A1(n2788), .A2(read_address_1[2]), .ZN(n1915) );
  AND2_X1 U1729 ( .A1(n2789), .A2(read_address_1[2]), .ZN(n1914) );
  AND2_X1 U1730 ( .A1(n2793), .A2(read_address_1[2]), .ZN(n1920) );
  INV_X1 U1731 ( .A(n1620), .ZN(n1616) );
  AOI22_X1 U1732 ( .A1(n2947), .A2(\bank_register[30][16] ), .B1(n2958), .B2(
        \bank_register[22][16] ), .ZN(n1620) );
  INV_X1 U1733 ( .A(n1583), .ZN(n1579) );
  AOI22_X1 U1734 ( .A1(n2947), .A2(\bank_register[30][17] ), .B1(n2958), .B2(
        \bank_register[22][17] ), .ZN(n1583) );
  INV_X1 U1735 ( .A(n1536), .ZN(n1532) );
  AOI22_X1 U1736 ( .A1(n2947), .A2(\bank_register[31][18] ), .B1(n2958), .B2(
        \bank_register[23][18] ), .ZN(n1536) );
  INV_X1 U1737 ( .A(n1509), .ZN(n1505) );
  AOI22_X1 U1738 ( .A1(n2947), .A2(\bank_register[30][19] ), .B1(n2958), .B2(
        \bank_register[22][19] ), .ZN(n1509) );
  INV_X1 U1739 ( .A(n1472), .ZN(n1468) );
  AOI22_X1 U1740 ( .A1(n2948), .A2(\bank_register[30][1] ), .B1(n2959), .B2(
        \bank_register[22][1] ), .ZN(n1472) );
  INV_X1 U1741 ( .A(n1462), .ZN(n1458) );
  AOI22_X1 U1742 ( .A1(n2948), .A2(\bank_register[31][1] ), .B1(n2959), .B2(
        \bank_register[23][1] ), .ZN(n1462) );
  INV_X1 U1743 ( .A(n1065), .ZN(n1061) );
  AOI22_X1 U1744 ( .A1(n2950), .A2(\bank_register[30][2] ), .B1(n2961), .B2(
        \bank_register[22][2] ), .ZN(n1065) );
  INV_X1 U1745 ( .A(n1055), .ZN(n1051) );
  AOI22_X1 U1746 ( .A1(n2950), .A2(\bank_register[31][2] ), .B1(n2961), .B2(
        \bank_register[23][2] ), .ZN(n1055) );
  INV_X1 U1747 ( .A(n1768), .ZN(n1764) );
  AOI22_X1 U1748 ( .A1(n2950), .A2(\bank_register[30][12] ), .B1(n2961), .B2(
        \bank_register[22][12] ), .ZN(n1768) );
  INV_X1 U1749 ( .A(n1721), .ZN(n1717) );
  AOI22_X1 U1750 ( .A1(n2949), .A2(\bank_register[31][13] ), .B1(n2960), .B2(
        \bank_register[23][13] ), .ZN(n1721) );
  INV_X1 U1751 ( .A(n1694), .ZN(n1690) );
  AOI22_X1 U1752 ( .A1(n2949), .A2(\bank_register[30][14] ), .B1(n2960), .B2(
        \bank_register[22][14] ), .ZN(n1694) );
  INV_X1 U1753 ( .A(n1684), .ZN(n1680) );
  AOI22_X1 U1754 ( .A1(n2949), .A2(\bank_register[31][14] ), .B1(n2961), .B2(
        \bank_register[23][14] ), .ZN(n1684) );
  INV_X1 U1755 ( .A(n1657), .ZN(n1653) );
  AOI22_X1 U1756 ( .A1(n2949), .A2(\bank_register[30][15] ), .B1(n2960), .B2(
        \bank_register[22][15] ), .ZN(n1657) );
  INV_X1 U1757 ( .A(n1647), .ZN(n1643) );
  AOI22_X1 U1758 ( .A1(n2948), .A2(\bank_register[31][15] ), .B1(n2959), .B2(
        \bank_register[23][15] ), .ZN(n1647) );
  INV_X1 U1759 ( .A(n1610), .ZN(n1606) );
  AOI22_X1 U1760 ( .A1(n2949), .A2(\bank_register[31][16] ), .B1(n2960), .B2(
        \bank_register[23][16] ), .ZN(n1610) );
  INV_X1 U1761 ( .A(n1573), .ZN(n1569) );
  AOI22_X1 U1762 ( .A1(n2948), .A2(\bank_register[31][17] ), .B1(n2959), .B2(
        \bank_register[23][17] ), .ZN(n1573) );
  INV_X1 U1763 ( .A(n1546), .ZN(n1542) );
  AOI22_X1 U1764 ( .A1(n2948), .A2(\bank_register[30][18] ), .B1(n2959), .B2(
        \bank_register[22][18] ), .ZN(n1546) );
  INV_X1 U1765 ( .A(n1499), .ZN(n1495) );
  AOI22_X1 U1766 ( .A1(n2948), .A2(\bank_register[31][19] ), .B1(n2959), .B2(
        \bank_register[23][19] ), .ZN(n1499) );
  INV_X1 U1767 ( .A(n1435), .ZN(n1431) );
  AOI22_X1 U1768 ( .A1(n2948), .A2(\bank_register[30][20] ), .B1(n2959), .B2(
        \bank_register[22][20] ), .ZN(n1435) );
  INV_X1 U1769 ( .A(n1425), .ZN(n1421) );
  AOI22_X1 U1770 ( .A1(n2948), .A2(\bank_register[31][20] ), .B1(n2959), .B2(
        \bank_register[23][20] ), .ZN(n1425) );
  INV_X1 U1771 ( .A(n1398), .ZN(n1394) );
  AOI22_X1 U1772 ( .A1(n2950), .A2(\bank_register[30][21] ), .B1(n2961), .B2(
        \bank_register[22][21] ), .ZN(n1398) );
  INV_X1 U1773 ( .A(n1388), .ZN(n1384) );
  AOI22_X1 U1774 ( .A1(n2948), .A2(\bank_register[31][21] ), .B1(n2959), .B2(
        \bank_register[23][21] ), .ZN(n1388) );
  INV_X1 U1775 ( .A(n1361), .ZN(n1357) );
  AOI22_X1 U1776 ( .A1(n2948), .A2(\bank_register[30][22] ), .B1(n2959), .B2(
        \bank_register[22][22] ), .ZN(n1361) );
  INV_X1 U1777 ( .A(n1351), .ZN(n1347) );
  AOI22_X1 U1778 ( .A1(n2948), .A2(\bank_register[31][22] ), .B1(n2959), .B2(
        \bank_register[23][22] ), .ZN(n1351) );
  INV_X1 U1779 ( .A(n1324), .ZN(n1320) );
  AOI22_X1 U1780 ( .A1(n2948), .A2(\bank_register[30][23] ), .B1(n2959), .B2(
        \bank_register[22][23] ), .ZN(n1324) );
  INV_X1 U1781 ( .A(n1314), .ZN(n1310) );
  AOI22_X1 U1782 ( .A1(n2948), .A2(\bank_register[31][23] ), .B1(n2960), .B2(
        \bank_register[23][23] ), .ZN(n1314) );
  INV_X1 U1783 ( .A(n1287), .ZN(n1283) );
  AOI22_X1 U1784 ( .A1(n2949), .A2(\bank_register[30][24] ), .B1(n2960), .B2(
        \bank_register[22][24] ), .ZN(n1287) );
  INV_X1 U1785 ( .A(n1277), .ZN(n1273) );
  AOI22_X1 U1786 ( .A1(n2949), .A2(\bank_register[31][24] ), .B1(n2960), .B2(
        \bank_register[23][24] ), .ZN(n1277) );
  INV_X1 U1787 ( .A(n1250), .ZN(n1246) );
  AOI22_X1 U1788 ( .A1(n2949), .A2(\bank_register[30][25] ), .B1(n2960), .B2(
        \bank_register[22][25] ), .ZN(n1250) );
  INV_X1 U1789 ( .A(n1240), .ZN(n1236) );
  AOI22_X1 U1790 ( .A1(n2949), .A2(\bank_register[31][25] ), .B1(n2960), .B2(
        \bank_register[23][25] ), .ZN(n1240) );
  INV_X1 U1791 ( .A(n1213), .ZN(n1209) );
  AOI22_X1 U1792 ( .A1(n2949), .A2(\bank_register[30][26] ), .B1(n2960), .B2(
        \bank_register[22][26] ), .ZN(n1213) );
  INV_X1 U1793 ( .A(n1203), .ZN(n1199) );
  AOI22_X1 U1794 ( .A1(n2949), .A2(\bank_register[31][26] ), .B1(n2960), .B2(
        \bank_register[23][26] ), .ZN(n1203) );
  INV_X1 U1795 ( .A(n1176), .ZN(n1172) );
  AOI22_X1 U1796 ( .A1(n2949), .A2(\bank_register[30][27] ), .B1(n2960), .B2(
        \bank_register[22][27] ), .ZN(n1176) );
  INV_X1 U1797 ( .A(n1166), .ZN(n1162) );
  AOI22_X1 U1798 ( .A1(n2949), .A2(\bank_register[31][27] ), .B1(n2961), .B2(
        \bank_register[23][27] ), .ZN(n1166) );
  INV_X1 U1799 ( .A(n1139), .ZN(n1135) );
  AOI22_X1 U1800 ( .A1(n2950), .A2(\bank_register[30][28] ), .B1(n2961), .B2(
        \bank_register[22][28] ), .ZN(n1139) );
  INV_X1 U1801 ( .A(n1129), .ZN(n1125) );
  AOI22_X1 U1802 ( .A1(n2950), .A2(\bank_register[31][28] ), .B1(n2961), .B2(
        \bank_register[23][28] ), .ZN(n1129) );
  INV_X1 U1803 ( .A(n1102), .ZN(n1098) );
  AOI22_X1 U1804 ( .A1(n2950), .A2(\bank_register[30][29] ), .B1(n2961), .B2(
        \bank_register[22][29] ), .ZN(n1102) );
  INV_X1 U1805 ( .A(n1092), .ZN(n1088) );
  AOI22_X1 U1806 ( .A1(n2950), .A2(\bank_register[31][29] ), .B1(n2961), .B2(
        \bank_register[23][29] ), .ZN(n1092) );
  INV_X1 U1807 ( .A(n1028), .ZN(n1024) );
  AOI22_X1 U1808 ( .A1(n2950), .A2(\bank_register[30][30] ), .B1(n2961), .B2(
        \bank_register[22][30] ), .ZN(n1028) );
  INV_X1 U1809 ( .A(n1018), .ZN(n1014) );
  AOI22_X1 U1810 ( .A1(n2950), .A2(\bank_register[31][30] ), .B1(n2961), .B2(
        \bank_register[23][30] ), .ZN(n1018) );
  INV_X1 U1811 ( .A(n954), .ZN(n950) );
  AOI22_X1 U1812 ( .A1(n2951), .A2(\bank_register[30][3] ), .B1(n2962), .B2(
        \bank_register[22][3] ), .ZN(n954) );
  INV_X1 U1813 ( .A(n944), .ZN(n940) );
  AOI22_X1 U1814 ( .A1(n2951), .A2(\bank_register[31][3] ), .B1(n2962), .B2(
        \bank_register[23][3] ), .ZN(n944) );
  INV_X1 U1815 ( .A(n917), .ZN(n913) );
  AOI22_X1 U1816 ( .A1(n2951), .A2(\bank_register[30][4] ), .B1(n2962), .B2(
        \bank_register[22][4] ), .ZN(n917) );
  INV_X1 U1817 ( .A(n907), .ZN(n903) );
  AOI22_X1 U1818 ( .A1(n2951), .A2(\bank_register[31][4] ), .B1(n2962), .B2(
        \bank_register[23][4] ), .ZN(n907) );
  INV_X1 U1819 ( .A(n880), .ZN(n876) );
  AOI22_X1 U1820 ( .A1(n2951), .A2(\bank_register[30][5] ), .B1(n2962), .B2(
        \bank_register[22][5] ), .ZN(n880) );
  INV_X1 U1821 ( .A(n870), .ZN(n866) );
  AOI22_X1 U1822 ( .A1(n2951), .A2(\bank_register[31][5] ), .B1(n2962), .B2(
        \bank_register[23][5] ), .ZN(n870) );
  INV_X1 U1823 ( .A(n843), .ZN(n839) );
  AOI22_X1 U1824 ( .A1(n2951), .A2(\bank_register[30][6] ), .B1(n2963), .B2(
        \bank_register[22][6] ), .ZN(n843) );
  INV_X1 U1825 ( .A(n833), .ZN(n829) );
  AOI22_X1 U1826 ( .A1(n2951), .A2(\bank_register[31][6] ), .B1(n2963), .B2(
        \bank_register[23][6] ), .ZN(n833) );
  INV_X1 U1827 ( .A(n806), .ZN(n802) );
  AOI22_X1 U1828 ( .A1(n2951), .A2(\bank_register[30][7] ), .B1(n2963), .B2(
        \bank_register[22][7] ), .ZN(n806) );
  INV_X1 U1829 ( .A(n1842), .ZN(n1838) );
  AOI22_X1 U1830 ( .A1(n2951), .A2(\bank_register[30][10] ), .B1(n2963), .B2(
        \bank_register[22][10] ), .ZN(n1842) );
  INV_X1 U1831 ( .A(n1805), .ZN(n1801) );
  AOI22_X1 U1832 ( .A1(n2951), .A2(\bank_register[30][11] ), .B1(n2962), .B2(
        \bank_register[22][11] ), .ZN(n1805) );
  INV_X1 U1833 ( .A(n1795), .ZN(n1791) );
  AOI22_X1 U1834 ( .A1(n2951), .A2(\bank_register[31][11] ), .B1(n2962), .B2(
        \bank_register[23][11] ), .ZN(n1795) );
  INV_X1 U1835 ( .A(n1758), .ZN(n1754) );
  AOI22_X1 U1836 ( .A1(n2951), .A2(\bank_register[31][12] ), .B1(n2962), .B2(
        \bank_register[23][12] ), .ZN(n1758) );
  INV_X1 U1837 ( .A(n1731), .ZN(n1727) );
  AOI22_X1 U1838 ( .A1(n2950), .A2(\bank_register[30][13] ), .B1(n2962), .B2(
        \bank_register[22][13] ), .ZN(n1731) );
  INV_X1 U1839 ( .A(n991), .ZN(n987) );
  AOI22_X1 U1840 ( .A1(n2950), .A2(\bank_register[30][31] ), .B1(n2962), .B2(
        \bank_register[22][31] ), .ZN(n991) );
  INV_X1 U1841 ( .A(n981), .ZN(n977) );
  AOI22_X1 U1842 ( .A1(n2950), .A2(\bank_register[31][31] ), .B1(n2962), .B2(
        \bank_register[23][31] ), .ZN(n981) );
  INV_X1 U1843 ( .A(n1621), .ZN(n1615) );
  AOI22_X1 U1844 ( .A1(n2991), .A2(\bank_register[14][16] ), .B1(n3002), .B2(
        \bank_register[26][16] ), .ZN(n1621) );
  INV_X1 U1845 ( .A(n1584), .ZN(n1578) );
  AOI22_X1 U1846 ( .A1(n2991), .A2(\bank_register[14][17] ), .B1(n3002), .B2(
        \bank_register[26][17] ), .ZN(n1584) );
  INV_X1 U1847 ( .A(n1537), .ZN(n1531) );
  AOI22_X1 U1848 ( .A1(n2991), .A2(\bank_register[15][18] ), .B1(n3002), .B2(
        \bank_register[27][18] ), .ZN(n1537) );
  INV_X1 U1849 ( .A(n1510), .ZN(n1504) );
  AOI22_X1 U1850 ( .A1(n2991), .A2(\bank_register[14][19] ), .B1(n3002), .B2(
        \bank_register[26][19] ), .ZN(n1510) );
  INV_X1 U1851 ( .A(n1473), .ZN(n1467) );
  AOI22_X1 U1852 ( .A1(n2992), .A2(\bank_register[14][1] ), .B1(n3003), .B2(
        \bank_register[26][1] ), .ZN(n1473) );
  INV_X1 U1853 ( .A(n1463), .ZN(n1457) );
  AOI22_X1 U1854 ( .A1(n2992), .A2(\bank_register[15][1] ), .B1(n3003), .B2(
        \bank_register[27][1] ), .ZN(n1463) );
  INV_X1 U1855 ( .A(n1066), .ZN(n1060) );
  AOI22_X1 U1856 ( .A1(n2994), .A2(\bank_register[14][2] ), .B1(n3005), .B2(
        \bank_register[26][2] ), .ZN(n1066) );
  INV_X1 U1857 ( .A(n1056), .ZN(n1050) );
  AOI22_X1 U1858 ( .A1(n2994), .A2(\bank_register[15][2] ), .B1(n3005), .B2(
        \bank_register[27][2] ), .ZN(n1056) );
  INV_X1 U1859 ( .A(n1769), .ZN(n1763) );
  AOI22_X1 U1860 ( .A1(n2994), .A2(\bank_register[14][12] ), .B1(n3005), .B2(
        \bank_register[26][12] ), .ZN(n1769) );
  INV_X1 U1861 ( .A(n1722), .ZN(n1716) );
  AOI22_X1 U1862 ( .A1(n2993), .A2(\bank_register[15][13] ), .B1(n3004), .B2(
        \bank_register[27][13] ), .ZN(n1722) );
  INV_X1 U1863 ( .A(n1695), .ZN(n1689) );
  AOI22_X1 U1864 ( .A1(n2993), .A2(\bank_register[14][14] ), .B1(n3004), .B2(
        \bank_register[26][14] ), .ZN(n1695) );
  INV_X1 U1865 ( .A(n1685), .ZN(n1679) );
  AOI22_X1 U1866 ( .A1(n2993), .A2(\bank_register[15][14] ), .B1(n3005), .B2(
        \bank_register[27][14] ), .ZN(n1685) );
  INV_X1 U1867 ( .A(n1658), .ZN(n1652) );
  AOI22_X1 U1868 ( .A1(n2993), .A2(\bank_register[14][15] ), .B1(n3004), .B2(
        \bank_register[26][15] ), .ZN(n1658) );
  INV_X1 U1869 ( .A(n1648), .ZN(n1642) );
  AOI22_X1 U1870 ( .A1(n2992), .A2(\bank_register[15][15] ), .B1(n3003), .B2(
        \bank_register[27][15] ), .ZN(n1648) );
  INV_X1 U1871 ( .A(n1611), .ZN(n1605) );
  AOI22_X1 U1872 ( .A1(n2993), .A2(\bank_register[15][16] ), .B1(n3004), .B2(
        \bank_register[27][16] ), .ZN(n1611) );
  INV_X1 U1873 ( .A(n1574), .ZN(n1568) );
  AOI22_X1 U1874 ( .A1(n2992), .A2(\bank_register[15][17] ), .B1(n3003), .B2(
        \bank_register[27][17] ), .ZN(n1574) );
  INV_X1 U1875 ( .A(n1547), .ZN(n1541) );
  AOI22_X1 U1876 ( .A1(n2992), .A2(\bank_register[14][18] ), .B1(n3003), .B2(
        \bank_register[26][18] ), .ZN(n1547) );
  INV_X1 U1877 ( .A(n1500), .ZN(n1494) );
  AOI22_X1 U1878 ( .A1(n2992), .A2(\bank_register[15][19] ), .B1(n3003), .B2(
        \bank_register[27][19] ), .ZN(n1500) );
  INV_X1 U1879 ( .A(n1436), .ZN(n1430) );
  AOI22_X1 U1880 ( .A1(n2992), .A2(\bank_register[14][20] ), .B1(n3003), .B2(
        \bank_register[26][20] ), .ZN(n1436) );
  INV_X1 U1881 ( .A(n1426), .ZN(n1420) );
  AOI22_X1 U1882 ( .A1(n2992), .A2(\bank_register[15][20] ), .B1(n3003), .B2(
        \bank_register[27][20] ), .ZN(n1426) );
  INV_X1 U1883 ( .A(n1399), .ZN(n1393) );
  AOI22_X1 U1884 ( .A1(n2994), .A2(\bank_register[14][21] ), .B1(n3005), .B2(
        \bank_register[26][21] ), .ZN(n1399) );
  INV_X1 U1885 ( .A(n1389), .ZN(n1383) );
  AOI22_X1 U1886 ( .A1(n2992), .A2(\bank_register[15][21] ), .B1(n3003), .B2(
        \bank_register[27][21] ), .ZN(n1389) );
  INV_X1 U1887 ( .A(n1362), .ZN(n1356) );
  AOI22_X1 U1888 ( .A1(n2992), .A2(\bank_register[14][22] ), .B1(n3003), .B2(
        \bank_register[26][22] ), .ZN(n1362) );
  INV_X1 U1889 ( .A(n1352), .ZN(n1346) );
  AOI22_X1 U1890 ( .A1(n2992), .A2(\bank_register[15][22] ), .B1(n3003), .B2(
        \bank_register[27][22] ), .ZN(n1352) );
  INV_X1 U1891 ( .A(n1325), .ZN(n1319) );
  AOI22_X1 U1892 ( .A1(n2992), .A2(\bank_register[14][23] ), .B1(n3003), .B2(
        \bank_register[26][23] ), .ZN(n1325) );
  INV_X1 U1893 ( .A(n1315), .ZN(n1309) );
  AOI22_X1 U1894 ( .A1(n2992), .A2(\bank_register[15][23] ), .B1(n3004), .B2(
        \bank_register[27][23] ), .ZN(n1315) );
  INV_X1 U1895 ( .A(n1288), .ZN(n1282) );
  AOI22_X1 U1896 ( .A1(n2993), .A2(\bank_register[14][24] ), .B1(n3004), .B2(
        \bank_register[26][24] ), .ZN(n1288) );
  INV_X1 U1897 ( .A(n1278), .ZN(n1272) );
  AOI22_X1 U1898 ( .A1(n2993), .A2(\bank_register[15][24] ), .B1(n3004), .B2(
        \bank_register[27][24] ), .ZN(n1278) );
  INV_X1 U1899 ( .A(n1251), .ZN(n1245) );
  AOI22_X1 U1900 ( .A1(n2993), .A2(\bank_register[14][25] ), .B1(n3004), .B2(
        \bank_register[26][25] ), .ZN(n1251) );
  INV_X1 U1901 ( .A(n1241), .ZN(n1235) );
  AOI22_X1 U1902 ( .A1(n2993), .A2(\bank_register[15][25] ), .B1(n3004), .B2(
        \bank_register[27][25] ), .ZN(n1241) );
  INV_X1 U1903 ( .A(n1214), .ZN(n1208) );
  AOI22_X1 U1904 ( .A1(n2993), .A2(\bank_register[14][26] ), .B1(n3004), .B2(
        \bank_register[26][26] ), .ZN(n1214) );
  INV_X1 U1905 ( .A(n1204), .ZN(n1198) );
  AOI22_X1 U1906 ( .A1(n2993), .A2(\bank_register[15][26] ), .B1(n3004), .B2(
        \bank_register[27][26] ), .ZN(n1204) );
  INV_X1 U1907 ( .A(n1177), .ZN(n1171) );
  AOI22_X1 U1908 ( .A1(n2993), .A2(\bank_register[14][27] ), .B1(n3004), .B2(
        \bank_register[26][27] ), .ZN(n1177) );
  INV_X1 U1909 ( .A(n1167), .ZN(n1161) );
  AOI22_X1 U1910 ( .A1(n2993), .A2(\bank_register[15][27] ), .B1(n3005), .B2(
        \bank_register[27][27] ), .ZN(n1167) );
  INV_X1 U1911 ( .A(n1140), .ZN(n1134) );
  AOI22_X1 U1912 ( .A1(n2994), .A2(\bank_register[14][28] ), .B1(n3005), .B2(
        \bank_register[26][28] ), .ZN(n1140) );
  INV_X1 U1913 ( .A(n1130), .ZN(n1124) );
  AOI22_X1 U1914 ( .A1(n2994), .A2(\bank_register[15][28] ), .B1(n3005), .B2(
        \bank_register[27][28] ), .ZN(n1130) );
  INV_X1 U1915 ( .A(n1103), .ZN(n1097) );
  AOI22_X1 U1916 ( .A1(n2994), .A2(\bank_register[14][29] ), .B1(n3005), .B2(
        \bank_register[26][29] ), .ZN(n1103) );
  INV_X1 U1917 ( .A(n1093), .ZN(n1087) );
  AOI22_X1 U1918 ( .A1(n2994), .A2(\bank_register[15][29] ), .B1(n3005), .B2(
        \bank_register[27][29] ), .ZN(n1093) );
  INV_X1 U1919 ( .A(n1029), .ZN(n1023) );
  AOI22_X1 U1920 ( .A1(n2994), .A2(\bank_register[14][30] ), .B1(n3005), .B2(
        \bank_register[26][30] ), .ZN(n1029) );
  INV_X1 U1921 ( .A(n1019), .ZN(n1013) );
  AOI22_X1 U1922 ( .A1(n2994), .A2(\bank_register[15][30] ), .B1(n3005), .B2(
        \bank_register[27][30] ), .ZN(n1019) );
  INV_X1 U1923 ( .A(n955), .ZN(n949) );
  AOI22_X1 U1924 ( .A1(n2995), .A2(\bank_register[14][3] ), .B1(n3006), .B2(
        \bank_register[26][3] ), .ZN(n955) );
  INV_X1 U1925 ( .A(n945), .ZN(n939) );
  AOI22_X1 U1926 ( .A1(n2995), .A2(\bank_register[15][3] ), .B1(n3006), .B2(
        \bank_register[27][3] ), .ZN(n945) );
  INV_X1 U1927 ( .A(n918), .ZN(n912) );
  AOI22_X1 U1928 ( .A1(n2995), .A2(\bank_register[14][4] ), .B1(n3006), .B2(
        \bank_register[26][4] ), .ZN(n918) );
  INV_X1 U1929 ( .A(n908), .ZN(n902) );
  AOI22_X1 U1930 ( .A1(n2995), .A2(\bank_register[15][4] ), .B1(n3006), .B2(
        \bank_register[27][4] ), .ZN(n908) );
  INV_X1 U1931 ( .A(n881), .ZN(n875) );
  AOI22_X1 U1932 ( .A1(n2995), .A2(\bank_register[14][5] ), .B1(n3006), .B2(
        \bank_register[26][5] ), .ZN(n881) );
  INV_X1 U1933 ( .A(n871), .ZN(n865) );
  AOI22_X1 U1934 ( .A1(n2995), .A2(\bank_register[15][5] ), .B1(n3006), .B2(
        \bank_register[27][5] ), .ZN(n871) );
  INV_X1 U1935 ( .A(n844), .ZN(n838) );
  AOI22_X1 U1936 ( .A1(n2995), .A2(\bank_register[14][6] ), .B1(n3007), .B2(
        \bank_register[26][6] ), .ZN(n844) );
  INV_X1 U1937 ( .A(n834), .ZN(n828) );
  AOI22_X1 U1938 ( .A1(n2995), .A2(\bank_register[15][6] ), .B1(n3007), .B2(
        \bank_register[27][6] ), .ZN(n834) );
  INV_X1 U1939 ( .A(n807), .ZN(n801) );
  AOI22_X1 U1940 ( .A1(n2995), .A2(\bank_register[14][7] ), .B1(n3007), .B2(
        \bank_register[26][7] ), .ZN(n807) );
  INV_X1 U1941 ( .A(n1843), .ZN(n1837) );
  AOI22_X1 U1942 ( .A1(n2995), .A2(\bank_register[14][10] ), .B1(n3007), .B2(
        \bank_register[26][10] ), .ZN(n1843) );
  INV_X1 U1943 ( .A(n1806), .ZN(n1800) );
  AOI22_X1 U1944 ( .A1(n2995), .A2(\bank_register[14][11] ), .B1(n3006), .B2(
        \bank_register[26][11] ), .ZN(n1806) );
  INV_X1 U1945 ( .A(n1796), .ZN(n1790) );
  AOI22_X1 U1946 ( .A1(n2995), .A2(\bank_register[15][11] ), .B1(n3006), .B2(
        \bank_register[27][11] ), .ZN(n1796) );
  INV_X1 U1947 ( .A(n1759), .ZN(n1753) );
  AOI22_X1 U1948 ( .A1(n2995), .A2(\bank_register[15][12] ), .B1(n3006), .B2(
        \bank_register[27][12] ), .ZN(n1759) );
  INV_X1 U1949 ( .A(n1732), .ZN(n1726) );
  AOI22_X1 U1950 ( .A1(n2994), .A2(\bank_register[14][13] ), .B1(n3006), .B2(
        \bank_register[26][13] ), .ZN(n1732) );
  INV_X1 U1951 ( .A(n992), .ZN(n986) );
  AOI22_X1 U1952 ( .A1(n2994), .A2(\bank_register[14][31] ), .B1(n3006), .B2(
        \bank_register[26][31] ), .ZN(n992) );
  INV_X1 U1953 ( .A(n982), .ZN(n976) );
  AOI22_X1 U1954 ( .A1(n2994), .A2(\bank_register[15][31] ), .B1(n3006), .B2(
        \bank_register[27][31] ), .ZN(n982) );
  NAND4_X1 U1955 ( .A1(n2760), .A2(n2761), .A3(n2762), .A4(n2763), .ZN(
        data_reg_1[0]) );
  NAND2_X1 U1956 ( .A1(n2917), .A2(write_data[0]), .ZN(n2760) );
  OAI21_X1 U1957 ( .B1(n2770), .B2(n2771), .A(n2823), .ZN(n2762) );
  NAND4_X1 U1958 ( .A1(n2485), .A2(n2486), .A3(n2487), .A4(n2488), .ZN(
        data_reg_1[1]) );
  NAND2_X1 U1959 ( .A1(n2918), .A2(write_data[1]), .ZN(n2485) );
  OAI21_X1 U1960 ( .B1(n2493), .B2(n2494), .A(n2823), .ZN(n2487) );
  NAND4_X1 U1961 ( .A1(n2710), .A2(n2711), .A3(n2712), .A4(n2713), .ZN(
        data_reg_1[11]) );
  NAND2_X1 U1962 ( .A1(n2919), .A2(write_data[11]), .ZN(n2710) );
  OAI21_X1 U1963 ( .B1(n2718), .B2(n2719), .A(n2823), .ZN(n2712) );
  NAND4_X1 U1964 ( .A1(n2685), .A2(n2686), .A3(n2687), .A4(n2688), .ZN(
        data_reg_1[12]) );
  NAND2_X1 U1965 ( .A1(n2919), .A2(write_data[12]), .ZN(n2685) );
  OAI21_X1 U1966 ( .B1(n2693), .B2(n2694), .A(n2823), .ZN(n2687) );
  NAND4_X1 U1967 ( .A1(n2660), .A2(n2661), .A3(n2662), .A4(n2663), .ZN(
        data_reg_1[13]) );
  NAND2_X1 U1968 ( .A1(n2919), .A2(write_data[13]), .ZN(n2660) );
  OAI21_X1 U1969 ( .B1(n2668), .B2(n2669), .A(n2823), .ZN(n2662) );
  NAND4_X1 U1970 ( .A1(n2635), .A2(n2636), .A3(n2637), .A4(n2638), .ZN(
        data_reg_1[14]) );
  NAND2_X1 U1971 ( .A1(n2919), .A2(write_data[14]), .ZN(n2635) );
  OAI21_X1 U1972 ( .B1(n2643), .B2(n2644), .A(n2823), .ZN(n2637) );
  NAND4_X1 U1973 ( .A1(n2610), .A2(n2611), .A3(n2612), .A4(n2613), .ZN(
        data_reg_1[15]) );
  NAND2_X1 U1974 ( .A1(n2919), .A2(write_data[15]), .ZN(n2610) );
  OAI21_X1 U1975 ( .B1(n2618), .B2(n2619), .A(n2823), .ZN(n2612) );
  NAND4_X1 U1976 ( .A1(n2585), .A2(n2586), .A3(n2587), .A4(n2588), .ZN(
        data_reg_1[16]) );
  NAND2_X1 U1977 ( .A1(n2919), .A2(write_data[16]), .ZN(n2585) );
  OAI21_X1 U1978 ( .B1(n2593), .B2(n2594), .A(n2823), .ZN(n2587) );
  NAND4_X1 U1979 ( .A1(n2560), .A2(n2561), .A3(n2562), .A4(n2563), .ZN(
        data_reg_1[17]) );
  NAND2_X1 U1980 ( .A1(n2919), .A2(write_data[17]), .ZN(n2560) );
  OAI21_X1 U1981 ( .B1(n2568), .B2(n2569), .A(n2823), .ZN(n2562) );
  NAND4_X1 U1982 ( .A1(n2535), .A2(n2536), .A3(n2537), .A4(n2538), .ZN(
        data_reg_1[18]) );
  NAND2_X1 U1983 ( .A1(n2918), .A2(write_data[18]), .ZN(n2535) );
  OAI21_X1 U1984 ( .B1(n2543), .B2(n2544), .A(n2823), .ZN(n2537) );
  NAND4_X1 U1985 ( .A1(n2510), .A2(n2511), .A3(n2512), .A4(n2513), .ZN(
        data_reg_1[19]) );
  NAND2_X1 U1986 ( .A1(n2918), .A2(write_data[19]), .ZN(n2510) );
  OAI21_X1 U1987 ( .B1(n2518), .B2(n2519), .A(n2823), .ZN(n2512) );
  NAND4_X1 U1988 ( .A1(n2460), .A2(n2461), .A3(n2462), .A4(n2463), .ZN(
        data_reg_1[20]) );
  NAND2_X1 U1989 ( .A1(n2918), .A2(write_data[20]), .ZN(n2460) );
  OAI21_X1 U1990 ( .B1(n2468), .B2(n2469), .A(n2824), .ZN(n2462) );
  NAND4_X1 U1991 ( .A1(n2435), .A2(n2436), .A3(n2437), .A4(n2438), .ZN(
        data_reg_1[21]) );
  NAND2_X1 U1992 ( .A1(n2918), .A2(write_data[21]), .ZN(n2435) );
  OAI21_X1 U1993 ( .B1(n2443), .B2(n2444), .A(n2824), .ZN(n2437) );
  NAND4_X1 U1994 ( .A1(n2410), .A2(n2411), .A3(n2412), .A4(n2413), .ZN(
        data_reg_1[22]) );
  NAND2_X1 U1995 ( .A1(n2918), .A2(write_data[22]), .ZN(n2410) );
  OAI21_X1 U1996 ( .B1(n2418), .B2(n2419), .A(n2824), .ZN(n2412) );
  NAND4_X1 U1997 ( .A1(n2385), .A2(n2386), .A3(n2387), .A4(n2388), .ZN(
        data_reg_1[23]) );
  NAND2_X1 U1998 ( .A1(n2918), .A2(write_data[23]), .ZN(n2385) );
  OAI21_X1 U1999 ( .B1(n2393), .B2(n2394), .A(n2824), .ZN(n2387) );
  NAND4_X1 U2000 ( .A1(n2356), .A2(n2358), .A3(n2359), .A4(n2360), .ZN(
        data_reg_1[24]) );
  NAND2_X1 U2001 ( .A1(n2918), .A2(write_data[24]), .ZN(n2356) );
  OAI21_X1 U2002 ( .B1(n2367), .B2(n2368), .A(n2824), .ZN(n2359) );
  NAND4_X1 U2003 ( .A1(n2323), .A2(n2324), .A3(n2326), .A4(n2327), .ZN(
        data_reg_1[25]) );
  NAND2_X1 U2004 ( .A1(n2918), .A2(write_data[25]), .ZN(n2323) );
  OAI21_X1 U2005 ( .B1(n2334), .B2(n2335), .A(n2824), .ZN(n2326) );
  NAND4_X1 U2006 ( .A1(n2290), .A2(n2291), .A3(n2292), .A4(n2294), .ZN(
        data_reg_1[26]) );
  NAND2_X1 U2007 ( .A1(n2918), .A2(write_data[26]), .ZN(n2290) );
  OAI21_X1 U2008 ( .B1(n2300), .B2(n2302), .A(n2824), .ZN(n2292) );
  NAND4_X1 U2009 ( .A1(n2256), .A2(n2258), .A3(n2259), .A4(n2260), .ZN(
        data_reg_1[27]) );
  NAND2_X1 U2010 ( .A1(n2918), .A2(write_data[27]), .ZN(n2256) );
  OAI21_X1 U2011 ( .B1(n2267), .B2(n2268), .A(n2824), .ZN(n2259) );
  NAND4_X1 U2012 ( .A1(n2220), .A2(n2222), .A3(n2223), .A4(n2225), .ZN(
        data_reg_1[28]) );
  NAND2_X1 U2013 ( .A1(n2918), .A2(write_data[28]), .ZN(n2220) );
  OAI21_X1 U2014 ( .B1(n2232), .B2(n2234), .A(n2824), .ZN(n2223) );
  NAND4_X1 U2015 ( .A1(n2183), .A2(n2184), .A3(n2186), .A4(n2187), .ZN(
        data_reg_1[29]) );
  NAND2_X1 U2016 ( .A1(n2917), .A2(write_data[29]), .ZN(n2183) );
  OAI21_X1 U2017 ( .B1(n2195), .B2(n2196), .A(n2824), .ZN(n2186) );
  NAND4_X1 U2018 ( .A1(n2122), .A2(n2123), .A3(n2124), .A4(n2125), .ZN(
        data_reg_1[30]) );
  NAND2_X1 U2019 ( .A1(n2917), .A2(write_data[30]), .ZN(n2122) );
  OAI21_X1 U2020 ( .B1(n2130), .B2(n2131), .A(n2824), .ZN(n2124) );
  NAND4_X1 U2021 ( .A1(n2097), .A2(n2098), .A3(n2099), .A4(n2100), .ZN(
        data_reg_1[31]) );
  NAND2_X1 U2022 ( .A1(n2918), .A2(write_data[31]), .ZN(n2097) );
  OAI21_X1 U2023 ( .B1(n2105), .B2(n2106), .A(n2825), .ZN(n2099) );
  NAND4_X1 U2024 ( .A1(n2147), .A2(n2148), .A3(n2149), .A4(n2150), .ZN(
        data_reg_1[2]) );
  NAND2_X1 U2025 ( .A1(n2917), .A2(write_data[2]), .ZN(n2147) );
  OAI21_X1 U2026 ( .B1(n2157), .B2(n2159), .A(n2824), .ZN(n2149) );
  NAND4_X1 U2027 ( .A1(n2072), .A2(n2073), .A3(n2074), .A4(n2075), .ZN(
        data_reg_1[3]) );
  NAND2_X1 U2028 ( .A1(n2917), .A2(write_data[3]), .ZN(n2072) );
  OAI21_X1 U2029 ( .B1(n2080), .B2(n2081), .A(n2825), .ZN(n2074) );
  NAND4_X1 U2030 ( .A1(n2047), .A2(n2048), .A3(n2049), .A4(n2050), .ZN(
        data_reg_1[4]) );
  NAND2_X1 U2031 ( .A1(n2917), .A2(write_data[4]), .ZN(n2047) );
  OAI21_X1 U2032 ( .B1(n2055), .B2(n2056), .A(n2825), .ZN(n2049) );
  NAND4_X1 U2033 ( .A1(n2022), .A2(n2023), .A3(n2024), .A4(n2025), .ZN(
        data_reg_1[5]) );
  NAND2_X1 U2034 ( .A1(n2917), .A2(write_data[5]), .ZN(n2022) );
  OAI21_X1 U2035 ( .B1(n2030), .B2(n2031), .A(n2825), .ZN(n2024) );
  NAND4_X1 U2036 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(
        data_reg_1[6]) );
  NAND2_X1 U2037 ( .A1(n2917), .A2(write_data[6]), .ZN(n1997) );
  OAI21_X1 U2038 ( .B1(n2005), .B2(n2006), .A(n2825), .ZN(n1999) );
  NAND4_X1 U2039 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .ZN(
        data_reg_1[7]) );
  NAND2_X1 U2040 ( .A1(n2917), .A2(write_data[7]), .ZN(n1972) );
  OAI21_X1 U2041 ( .B1(n1980), .B2(n1981), .A(n2825), .ZN(n1974) );
  NAND4_X1 U2042 ( .A1(n1947), .A2(n1948), .A3(n1949), .A4(n1950), .ZN(
        data_reg_1[8]) );
  NAND2_X1 U2043 ( .A1(n2917), .A2(write_data[8]), .ZN(n1947) );
  OAI21_X1 U2044 ( .B1(n1955), .B2(n1956), .A(n2825), .ZN(n1949) );
  NAND4_X1 U2045 ( .A1(n1904), .A2(n1905), .A3(n1906), .A4(n1907), .ZN(
        data_reg_1[9]) );
  NAND2_X1 U2046 ( .A1(n2917), .A2(write_data[9]), .ZN(n1904) );
  OAI21_X1 U2047 ( .B1(n1921), .B2(n1922), .A(n2825), .ZN(n1906) );
  NAND4_X1 U2048 ( .A1(n2735), .A2(n2736), .A3(n2737), .A4(n2738), .ZN(
        data_reg_1[10]) );
  NAND2_X1 U2049 ( .A1(n2919), .A2(write_data[10]), .ZN(n2735) );
  OAI21_X1 U2050 ( .B1(n2743), .B2(n2744), .A(n2823), .ZN(n2737) );
  INV_X1 U2051 ( .A(write_address[0]), .ZN(n678) );
  INV_X1 U2052 ( .A(write_address[1]), .ZN(n676) );
  INV_X1 U2053 ( .A(write_address[2]), .ZN(n677) );
  INV_X1 U2054 ( .A(\bank_register[2][0] ), .ZN(n1894) );
  INV_X1 U2055 ( .A(\bank_register[10][0] ), .ZN(n1903) );
  INV_X1 U2056 ( .A(\bank_register[3][0] ), .ZN(n1873) );
  INV_X1 U2057 ( .A(\bank_register[11][0] ), .ZN(n1877) );
  INV_X1 U2058 ( .A(\bank_register[2][1] ), .ZN(n1471) );
  INV_X1 U2059 ( .A(\bank_register[10][1] ), .ZN(n1475) );
  INV_X1 U2060 ( .A(\bank_register[3][1] ), .ZN(n1461) );
  INV_X1 U2061 ( .A(\bank_register[11][1] ), .ZN(n1465) );
  INV_X1 U2062 ( .A(\bank_register[2][2] ), .ZN(n1064) );
  INV_X1 U2063 ( .A(\bank_register[10][2] ), .ZN(n1068) );
  INV_X1 U2064 ( .A(\bank_register[3][2] ), .ZN(n1054) );
  INV_X1 U2065 ( .A(\bank_register[11][2] ), .ZN(n1058) );
  INV_X1 U2066 ( .A(\bank_register[2][3] ), .ZN(n953) );
  INV_X1 U2067 ( .A(\bank_register[10][3] ), .ZN(n957) );
  INV_X1 U2068 ( .A(\bank_register[3][3] ), .ZN(n943) );
  INV_X1 U2069 ( .A(\bank_register[11][3] ), .ZN(n947) );
  INV_X1 U2070 ( .A(\bank_register[2][4] ), .ZN(n916) );
  INV_X1 U2071 ( .A(\bank_register[10][4] ), .ZN(n920) );
  INV_X1 U2072 ( .A(\bank_register[3][4] ), .ZN(n906) );
  INV_X1 U2073 ( .A(\bank_register[11][4] ), .ZN(n910) );
  INV_X1 U2074 ( .A(\bank_register[2][5] ), .ZN(n879) );
  INV_X1 U2075 ( .A(\bank_register[10][5] ), .ZN(n883) );
  INV_X1 U2076 ( .A(\bank_register[3][5] ), .ZN(n869) );
  INV_X1 U2077 ( .A(\bank_register[11][5] ), .ZN(n873) );
  INV_X1 U2078 ( .A(\bank_register[2][6] ), .ZN(n842) );
  INV_X1 U2079 ( .A(\bank_register[10][6] ), .ZN(n846) );
  INV_X1 U2080 ( .A(\bank_register[3][6] ), .ZN(n832) );
  INV_X1 U2081 ( .A(\bank_register[11][6] ), .ZN(n836) );
  INV_X1 U2082 ( .A(\bank_register[2][7] ), .ZN(n805) );
  INV_X1 U2083 ( .A(\bank_register[10][7] ), .ZN(n809) );
  INV_X1 U2084 ( .A(\bank_register[3][7] ), .ZN(n795) );
  INV_X1 U2085 ( .A(\bank_register[11][7] ), .ZN(n799) );
  INV_X1 U2086 ( .A(\bank_register[2][8] ), .ZN(n768) );
  INV_X1 U2087 ( .A(\bank_register[10][8] ), .ZN(n772) );
  INV_X1 U2088 ( .A(\bank_register[3][8] ), .ZN(n758) );
  INV_X1 U2089 ( .A(\bank_register[11][8] ), .ZN(n762) );
  INV_X1 U2090 ( .A(\bank_register[2][9] ), .ZN(n731) );
  INV_X1 U2091 ( .A(\bank_register[10][9] ), .ZN(n735) );
  INV_X1 U2092 ( .A(\bank_register[3][9] ), .ZN(n721) );
  INV_X1 U2093 ( .A(\bank_register[11][9] ), .ZN(n725) );
  INV_X1 U2094 ( .A(\bank_register[2][10] ), .ZN(n1841) );
  INV_X1 U2095 ( .A(\bank_register[10][10] ), .ZN(n1845) );
  INV_X1 U2096 ( .A(\bank_register[3][10] ), .ZN(n1831) );
  INV_X1 U2097 ( .A(\bank_register[11][10] ), .ZN(n1835) );
  INV_X1 U2098 ( .A(\bank_register[2][11] ), .ZN(n1804) );
  INV_X1 U2099 ( .A(\bank_register[10][11] ), .ZN(n1808) );
  INV_X1 U2100 ( .A(\bank_register[3][11] ), .ZN(n1794) );
  INV_X1 U2101 ( .A(\bank_register[11][11] ), .ZN(n1798) );
  INV_X1 U2102 ( .A(\bank_register[2][12] ), .ZN(n1767) );
  INV_X1 U2103 ( .A(\bank_register[10][12] ), .ZN(n1771) );
  INV_X1 U2104 ( .A(\bank_register[3][12] ), .ZN(n1757) );
  INV_X1 U2105 ( .A(\bank_register[11][12] ), .ZN(n1761) );
  INV_X1 U2106 ( .A(\bank_register[2][13] ), .ZN(n1730) );
  INV_X1 U2107 ( .A(\bank_register[10][13] ), .ZN(n1734) );
  INV_X1 U2108 ( .A(\bank_register[3][13] ), .ZN(n1720) );
  INV_X1 U2109 ( .A(\bank_register[11][13] ), .ZN(n1724) );
  INV_X1 U2110 ( .A(\bank_register[2][14] ), .ZN(n1693) );
  INV_X1 U2111 ( .A(\bank_register[10][14] ), .ZN(n1697) );
  INV_X1 U2112 ( .A(\bank_register[3][14] ), .ZN(n1683) );
  INV_X1 U2113 ( .A(\bank_register[11][14] ), .ZN(n1687) );
  INV_X1 U2114 ( .A(\bank_register[2][15] ), .ZN(n1656) );
  INV_X1 U2115 ( .A(\bank_register[10][15] ), .ZN(n1660) );
  INV_X1 U2116 ( .A(\bank_register[3][15] ), .ZN(n1646) );
  INV_X1 U2117 ( .A(\bank_register[11][15] ), .ZN(n1650) );
  INV_X1 U2118 ( .A(\bank_register[2][16] ), .ZN(n1619) );
  INV_X1 U2119 ( .A(\bank_register[10][16] ), .ZN(n1623) );
  INV_X1 U2120 ( .A(\bank_register[3][16] ), .ZN(n1609) );
  INV_X1 U2121 ( .A(\bank_register[11][16] ), .ZN(n1613) );
  INV_X1 U2122 ( .A(\bank_register[2][17] ), .ZN(n1582) );
  INV_X1 U2123 ( .A(\bank_register[10][17] ), .ZN(n1586) );
  INV_X1 U2124 ( .A(\bank_register[3][17] ), .ZN(n1572) );
  INV_X1 U2125 ( .A(\bank_register[11][17] ), .ZN(n1576) );
  INV_X1 U2126 ( .A(\bank_register[2][18] ), .ZN(n1545) );
  INV_X1 U2127 ( .A(\bank_register[10][18] ), .ZN(n1549) );
  INV_X1 U2128 ( .A(\bank_register[3][18] ), .ZN(n1535) );
  INV_X1 U2129 ( .A(\bank_register[11][18] ), .ZN(n1539) );
  INV_X1 U2130 ( .A(\bank_register[2][19] ), .ZN(n1508) );
  INV_X1 U2131 ( .A(\bank_register[10][19] ), .ZN(n1512) );
  INV_X1 U2132 ( .A(\bank_register[3][19] ), .ZN(n1498) );
  INV_X1 U2133 ( .A(\bank_register[11][19] ), .ZN(n1502) );
  INV_X1 U2134 ( .A(\bank_register[2][20] ), .ZN(n1434) );
  INV_X1 U2135 ( .A(\bank_register[10][20] ), .ZN(n1438) );
  INV_X1 U2136 ( .A(\bank_register[3][20] ), .ZN(n1424) );
  INV_X1 U2137 ( .A(\bank_register[11][20] ), .ZN(n1428) );
  INV_X1 U2138 ( .A(\bank_register[2][21] ), .ZN(n1397) );
  INV_X1 U2139 ( .A(\bank_register[10][21] ), .ZN(n1401) );
  INV_X1 U2140 ( .A(\bank_register[3][21] ), .ZN(n1387) );
  INV_X1 U2141 ( .A(\bank_register[11][21] ), .ZN(n1391) );
  INV_X1 U2142 ( .A(\bank_register[2][22] ), .ZN(n1360) );
  INV_X1 U2143 ( .A(\bank_register[10][22] ), .ZN(n1364) );
  INV_X1 U2144 ( .A(\bank_register[3][22] ), .ZN(n1350) );
  INV_X1 U2145 ( .A(\bank_register[11][22] ), .ZN(n1354) );
  INV_X1 U2146 ( .A(\bank_register[2][23] ), .ZN(n1323) );
  INV_X1 U2147 ( .A(\bank_register[10][23] ), .ZN(n1327) );
  INV_X1 U2148 ( .A(\bank_register[3][23] ), .ZN(n1313) );
  INV_X1 U2149 ( .A(\bank_register[11][23] ), .ZN(n1317) );
  INV_X1 U2150 ( .A(\bank_register[2][24] ), .ZN(n1286) );
  INV_X1 U2151 ( .A(\bank_register[10][24] ), .ZN(n1290) );
  INV_X1 U2152 ( .A(\bank_register[3][24] ), .ZN(n1276) );
  INV_X1 U2153 ( .A(\bank_register[11][24] ), .ZN(n1280) );
  INV_X1 U2154 ( .A(\bank_register[2][25] ), .ZN(n1249) );
  INV_X1 U2155 ( .A(\bank_register[10][25] ), .ZN(n1253) );
  INV_X1 U2156 ( .A(\bank_register[3][25] ), .ZN(n1239) );
  INV_X1 U2157 ( .A(\bank_register[11][25] ), .ZN(n1243) );
  INV_X1 U2158 ( .A(\bank_register[2][26] ), .ZN(n1212) );
  INV_X1 U2159 ( .A(\bank_register[10][26] ), .ZN(n1216) );
  INV_X1 U2160 ( .A(\bank_register[3][26] ), .ZN(n1202) );
  INV_X1 U2161 ( .A(\bank_register[11][26] ), .ZN(n1206) );
  INV_X1 U2162 ( .A(\bank_register[2][27] ), .ZN(n1175) );
  INV_X1 U2163 ( .A(\bank_register[10][27] ), .ZN(n1179) );
  INV_X1 U2164 ( .A(\bank_register[3][27] ), .ZN(n1165) );
  INV_X1 U2165 ( .A(\bank_register[11][27] ), .ZN(n1169) );
  INV_X1 U2166 ( .A(\bank_register[2][28] ), .ZN(n1138) );
  INV_X1 U2167 ( .A(\bank_register[10][28] ), .ZN(n1142) );
  INV_X1 U2168 ( .A(\bank_register[3][28] ), .ZN(n1128) );
  INV_X1 U2169 ( .A(\bank_register[11][28] ), .ZN(n1132) );
  INV_X1 U2170 ( .A(\bank_register[2][29] ), .ZN(n1101) );
  INV_X1 U2171 ( .A(\bank_register[10][29] ), .ZN(n1105) );
  INV_X1 U2172 ( .A(\bank_register[3][29] ), .ZN(n1091) );
  INV_X1 U2173 ( .A(\bank_register[11][29] ), .ZN(n1095) );
  INV_X1 U2174 ( .A(\bank_register[2][30] ), .ZN(n1027) );
  INV_X1 U2175 ( .A(\bank_register[10][30] ), .ZN(n1031) );
  INV_X1 U2176 ( .A(\bank_register[3][30] ), .ZN(n1017) );
  INV_X1 U2177 ( .A(\bank_register[11][30] ), .ZN(n1021) );
  INV_X1 U2178 ( .A(\bank_register[2][31] ), .ZN(n990) );
  INV_X1 U2205 ( .A(\bank_register[10][31] ), .ZN(n994) );
  INV_X1 U2206 ( .A(\bank_register[3][31] ), .ZN(n980) );
  INV_X1 U2207 ( .A(\bank_register[11][31] ), .ZN(n984) );
  INV_X1 U2208 ( .A(\bank_register[17][0] ), .ZN(n1862) );
  INV_X1 U2209 ( .A(\bank_register[5][0] ), .ZN(n1865) );
  INV_X1 U2210 ( .A(\bank_register[17][1] ), .ZN(n1451) );
  INV_X1 U2211 ( .A(\bank_register[5][1] ), .ZN(n1454) );
  INV_X1 U2212 ( .A(\bank_register[17][2] ), .ZN(n1044) );
  INV_X1 U2213 ( .A(\bank_register[5][2] ), .ZN(n1047) );
  INV_X1 U2214 ( .A(\bank_register[17][3] ), .ZN(n933) );
  INV_X1 U2215 ( .A(\bank_register[5][3] ), .ZN(n936) );
  INV_X1 U2216 ( .A(\bank_register[17][4] ), .ZN(n896) );
  INV_X1 U2217 ( .A(\bank_register[5][4] ), .ZN(n899) );
  INV_X1 U2218 ( .A(\bank_register[17][5] ), .ZN(n859) );
  INV_X1 U2219 ( .A(\bank_register[5][5] ), .ZN(n862) );
  INV_X1 U2220 ( .A(\bank_register[17][6] ), .ZN(n822) );
  INV_X1 U2221 ( .A(\bank_register[5][6] ), .ZN(n825) );
  INV_X1 U2222 ( .A(\bank_register[17][7] ), .ZN(n785) );
  INV_X1 U2223 ( .A(\bank_register[5][7] ), .ZN(n788) );
  INV_X1 U2224 ( .A(\bank_register[17][8] ), .ZN(n748) );
  INV_X1 U2225 ( .A(\bank_register[5][8] ), .ZN(n751) );
  INV_X1 U2226 ( .A(\bank_register[17][9] ), .ZN(n706) );
  INV_X1 U2227 ( .A(\bank_register[5][9] ), .ZN(n713) );
  INV_X1 U2228 ( .A(\bank_register[17][10] ), .ZN(n1821) );
  INV_X1 U2229 ( .A(\bank_register[5][10] ), .ZN(n1824) );
  INV_X1 U2230 ( .A(\bank_register[17][11] ), .ZN(n1784) );
  INV_X1 U2231 ( .A(\bank_register[5][11] ), .ZN(n1787) );
  INV_X1 U2232 ( .A(\bank_register[17][12] ), .ZN(n1747) );
  INV_X1 U2233 ( .A(\bank_register[5][12] ), .ZN(n1750) );
  INV_X1 U2234 ( .A(\bank_register[17][13] ), .ZN(n1710) );
  INV_X1 U2235 ( .A(\bank_register[5][13] ), .ZN(n1713) );
  INV_X1 U2236 ( .A(\bank_register[17][14] ), .ZN(n1673) );
  INV_X1 U2237 ( .A(\bank_register[5][14] ), .ZN(n1676) );
  INV_X1 U2238 ( .A(\bank_register[17][15] ), .ZN(n1636) );
  INV_X1 U2239 ( .A(\bank_register[5][15] ), .ZN(n1639) );
  INV_X1 U2240 ( .A(\bank_register[17][16] ), .ZN(n1599) );
  INV_X1 U2241 ( .A(\bank_register[5][16] ), .ZN(n1602) );
  INV_X1 U2242 ( .A(\bank_register[17][17] ), .ZN(n1562) );
  INV_X1 U2243 ( .A(\bank_register[5][17] ), .ZN(n1565) );
  INV_X1 U2244 ( .A(\bank_register[17][18] ), .ZN(n1525) );
  INV_X1 U2245 ( .A(\bank_register[5][18] ), .ZN(n1528) );
  INV_X1 U2246 ( .A(\bank_register[17][19] ), .ZN(n1488) );
  INV_X1 U2247 ( .A(\bank_register[5][19] ), .ZN(n1491) );
  INV_X1 U2248 ( .A(\bank_register[17][20] ), .ZN(n1414) );
  INV_X1 U2249 ( .A(\bank_register[5][20] ), .ZN(n1417) );
  INV_X1 U2250 ( .A(\bank_register[17][21] ), .ZN(n1377) );
  INV_X1 U2251 ( .A(\bank_register[5][21] ), .ZN(n1380) );
  INV_X1 U2252 ( .A(\bank_register[17][22] ), .ZN(n1340) );
  INV_X1 U2253 ( .A(\bank_register[5][22] ), .ZN(n1343) );
  INV_X1 U2254 ( .A(\bank_register[17][23] ), .ZN(n1303) );
  INV_X1 U2255 ( .A(\bank_register[5][23] ), .ZN(n1306) );
  INV_X1 U2256 ( .A(\bank_register[17][24] ), .ZN(n1266) );
  INV_X1 U2257 ( .A(\bank_register[5][24] ), .ZN(n1269) );
  INV_X1 U2258 ( .A(\bank_register[17][25] ), .ZN(n1229) );
  INV_X1 U2259 ( .A(\bank_register[5][25] ), .ZN(n1232) );
  INV_X1 U2260 ( .A(\bank_register[17][26] ), .ZN(n1192) );
  INV_X1 U2261 ( .A(\bank_register[5][26] ), .ZN(n1195) );
  INV_X1 U2262 ( .A(\bank_register[17][27] ), .ZN(n1155) );
  INV_X1 U2263 ( .A(\bank_register[5][27] ), .ZN(n1158) );
  INV_X1 U2264 ( .A(\bank_register[17][28] ), .ZN(n1118) );
  INV_X1 U2265 ( .A(\bank_register[5][28] ), .ZN(n1121) );
  INV_X1 U2266 ( .A(\bank_register[17][29] ), .ZN(n1081) );
  INV_X1 U2267 ( .A(\bank_register[5][29] ), .ZN(n1084) );
  INV_X1 U2268 ( .A(\bank_register[17][30] ), .ZN(n1007) );
  INV_X1 U2269 ( .A(\bank_register[5][30] ), .ZN(n1010) );
  INV_X1 U2270 ( .A(\bank_register[17][31] ), .ZN(n970) );
  INV_X1 U2271 ( .A(\bank_register[5][31] ), .ZN(n973) );
  INV_X1 U2272 ( .A(\bank_register[9][0] ), .ZN(n1863) );
  INV_X1 U2273 ( .A(\bank_register[1][0] ), .ZN(n1866) );
  INV_X1 U2274 ( .A(\bank_register[9][1] ), .ZN(n1452) );
  INV_X1 U2275 ( .A(\bank_register[1][1] ), .ZN(n1455) );
  INV_X1 U2276 ( .A(\bank_register[9][2] ), .ZN(n1045) );
  INV_X1 U2277 ( .A(\bank_register[1][2] ), .ZN(n1048) );
  INV_X1 U2278 ( .A(\bank_register[9][3] ), .ZN(n934) );
  INV_X1 U2279 ( .A(\bank_register[1][3] ), .ZN(n937) );
  INV_X1 U2280 ( .A(\bank_register[9][4] ), .ZN(n897) );
  INV_X1 U2281 ( .A(\bank_register[1][4] ), .ZN(n900) );
  INV_X1 U2282 ( .A(\bank_register[9][5] ), .ZN(n860) );
  INV_X1 U2283 ( .A(\bank_register[1][5] ), .ZN(n863) );
  INV_X1 U2284 ( .A(\bank_register[9][6] ), .ZN(n823) );
  INV_X1 U2285 ( .A(\bank_register[1][6] ), .ZN(n826) );
  INV_X1 U2286 ( .A(\bank_register[9][7] ), .ZN(n786) );
  INV_X1 U2287 ( .A(\bank_register[1][7] ), .ZN(n789) );
  INV_X1 U2288 ( .A(\bank_register[9][8] ), .ZN(n749) );
  INV_X1 U2289 ( .A(\bank_register[1][8] ), .ZN(n752) );
  INV_X1 U2290 ( .A(\bank_register[9][9] ), .ZN(n708) );
  INV_X1 U2291 ( .A(\bank_register[1][9] ), .ZN(n715) );
  INV_X1 U2292 ( .A(\bank_register[9][10] ), .ZN(n1822) );
  INV_X1 U2293 ( .A(\bank_register[1][10] ), .ZN(n1825) );
  INV_X1 U2294 ( .A(\bank_register[9][11] ), .ZN(n1785) );
  INV_X1 U2295 ( .A(\bank_register[1][11] ), .ZN(n1788) );
  INV_X1 U2296 ( .A(\bank_register[9][12] ), .ZN(n1748) );
  INV_X1 U2297 ( .A(\bank_register[1][12] ), .ZN(n1751) );
  INV_X1 U2298 ( .A(\bank_register[9][13] ), .ZN(n1711) );
  INV_X1 U2299 ( .A(\bank_register[1][13] ), .ZN(n1714) );
  INV_X1 U2300 ( .A(\bank_register[9][14] ), .ZN(n1674) );
  INV_X1 U2301 ( .A(\bank_register[1][14] ), .ZN(n1677) );
  INV_X1 U2302 ( .A(\bank_register[9][15] ), .ZN(n1637) );
  INV_X1 U2303 ( .A(\bank_register[1][15] ), .ZN(n1640) );
  INV_X1 U2304 ( .A(\bank_register[9][16] ), .ZN(n1600) );
  INV_X1 U2305 ( .A(\bank_register[1][16] ), .ZN(n1603) );
  INV_X1 U2306 ( .A(\bank_register[9][17] ), .ZN(n1563) );
  INV_X1 U2307 ( .A(\bank_register[1][17] ), .ZN(n1566) );
  INV_X1 U2308 ( .A(\bank_register[9][18] ), .ZN(n1526) );
  INV_X1 U2309 ( .A(\bank_register[1][18] ), .ZN(n1529) );
  INV_X1 U2310 ( .A(\bank_register[9][19] ), .ZN(n1489) );
  INV_X1 U2311 ( .A(\bank_register[1][19] ), .ZN(n1492) );
  INV_X1 U2312 ( .A(\bank_register[9][20] ), .ZN(n1415) );
  INV_X1 U2313 ( .A(\bank_register[1][20] ), .ZN(n1418) );
  INV_X1 U2314 ( .A(\bank_register[9][21] ), .ZN(n1378) );
  INV_X1 U2315 ( .A(\bank_register[1][21] ), .ZN(n1381) );
  INV_X1 U2316 ( .A(\bank_register[9][22] ), .ZN(n1341) );
  INV_X1 U2317 ( .A(\bank_register[1][22] ), .ZN(n1344) );
  INV_X1 U2318 ( .A(\bank_register[9][23] ), .ZN(n1304) );
  INV_X1 U2319 ( .A(\bank_register[1][23] ), .ZN(n1307) );
  INV_X1 U2320 ( .A(\bank_register[9][24] ), .ZN(n1267) );
  INV_X1 U2321 ( .A(\bank_register[1][24] ), .ZN(n1270) );
  INV_X1 U2322 ( .A(\bank_register[9][25] ), .ZN(n1230) );
  INV_X1 U2323 ( .A(\bank_register[1][25] ), .ZN(n1233) );
  INV_X1 U2324 ( .A(\bank_register[9][26] ), .ZN(n1193) );
  INV_X1 U2325 ( .A(\bank_register[1][26] ), .ZN(n1196) );
  INV_X1 U2326 ( .A(\bank_register[9][27] ), .ZN(n1156) );
  INV_X1 U2327 ( .A(\bank_register[1][27] ), .ZN(n1159) );
  INV_X1 U2328 ( .A(\bank_register[9][28] ), .ZN(n1119) );
  INV_X1 U2329 ( .A(\bank_register[1][28] ), .ZN(n1122) );
  INV_X1 U2330 ( .A(\bank_register[9][29] ), .ZN(n1082) );
  INV_X1 U2331 ( .A(\bank_register[1][29] ), .ZN(n1085) );
  INV_X1 U2332 ( .A(\bank_register[9][30] ), .ZN(n1008) );
  INV_X1 U2333 ( .A(\bank_register[1][30] ), .ZN(n1011) );
  INV_X1 U2334 ( .A(\bank_register[9][31] ), .ZN(n971) );
  INV_X1 U2335 ( .A(\bank_register[1][31] ), .ZN(n974) );
  INV_X1 U2336 ( .A(\bank_register[6][0] ), .ZN(n1893) );
  INV_X1 U2337 ( .A(\bank_register[18][0] ), .ZN(n1902) );
  INV_X1 U2338 ( .A(\bank_register[7][0] ), .ZN(n1872) );
  INV_X1 U2339 ( .A(\bank_register[19][0] ), .ZN(n1876) );
  INV_X1 U2340 ( .A(\bank_register[6][1] ), .ZN(n1470) );
  INV_X1 U2341 ( .A(\bank_register[18][1] ), .ZN(n1474) );
  INV_X1 U2342 ( .A(\bank_register[7][1] ), .ZN(n1460) );
  INV_X1 U2343 ( .A(\bank_register[19][1] ), .ZN(n1464) );
  INV_X1 U2344 ( .A(\bank_register[6][2] ), .ZN(n1063) );
  INV_X1 U2345 ( .A(\bank_register[18][2] ), .ZN(n1067) );
  INV_X1 U2346 ( .A(\bank_register[7][2] ), .ZN(n1053) );
  INV_X1 U2347 ( .A(\bank_register[19][2] ), .ZN(n1057) );
  INV_X1 U2348 ( .A(\bank_register[6][3] ), .ZN(n952) );
  INV_X1 U2349 ( .A(\bank_register[18][3] ), .ZN(n956) );
  INV_X1 U2350 ( .A(\bank_register[7][3] ), .ZN(n942) );
  INV_X1 U2351 ( .A(\bank_register[19][3] ), .ZN(n946) );
  INV_X1 U2352 ( .A(\bank_register[6][4] ), .ZN(n915) );
  INV_X1 U2353 ( .A(\bank_register[18][4] ), .ZN(n919) );
  INV_X1 U2354 ( .A(\bank_register[7][4] ), .ZN(n905) );
  INV_X1 U2355 ( .A(\bank_register[19][4] ), .ZN(n909) );
  INV_X1 U2356 ( .A(\bank_register[6][5] ), .ZN(n878) );
  INV_X1 U2357 ( .A(\bank_register[18][5] ), .ZN(n882) );
  INV_X1 U2358 ( .A(\bank_register[7][5] ), .ZN(n868) );
  INV_X1 U2359 ( .A(\bank_register[19][5] ), .ZN(n872) );
  INV_X1 U2360 ( .A(\bank_register[6][6] ), .ZN(n841) );
  INV_X1 U2361 ( .A(\bank_register[18][6] ), .ZN(n845) );
  INV_X1 U2362 ( .A(\bank_register[7][6] ), .ZN(n831) );
  INV_X1 U2363 ( .A(\bank_register[19][6] ), .ZN(n835) );
  INV_X1 U2364 ( .A(\bank_register[6][7] ), .ZN(n804) );
  INV_X1 U2365 ( .A(\bank_register[18][7] ), .ZN(n808) );
  INV_X1 U2366 ( .A(\bank_register[7][7] ), .ZN(n794) );
  INV_X1 U2367 ( .A(\bank_register[19][7] ), .ZN(n798) );
  INV_X1 U2368 ( .A(\bank_register[6][8] ), .ZN(n767) );
  INV_X1 U2369 ( .A(\bank_register[18][8] ), .ZN(n771) );
  INV_X1 U2370 ( .A(\bank_register[7][8] ), .ZN(n757) );
  INV_X1 U2371 ( .A(\bank_register[19][8] ), .ZN(n761) );
  INV_X1 U2372 ( .A(\bank_register[6][9] ), .ZN(n730) );
  INV_X1 U2373 ( .A(\bank_register[18][9] ), .ZN(n734) );
  INV_X1 U2374 ( .A(\bank_register[7][9] ), .ZN(n720) );
  INV_X1 U2375 ( .A(\bank_register[19][9] ), .ZN(n724) );
  INV_X1 U2376 ( .A(\bank_register[6][10] ), .ZN(n1840) );
  INV_X1 U2377 ( .A(\bank_register[18][10] ), .ZN(n1844) );
  INV_X1 U2378 ( .A(\bank_register[7][10] ), .ZN(n1830) );
  INV_X1 U2379 ( .A(\bank_register[19][10] ), .ZN(n1834) );
  INV_X1 U2380 ( .A(\bank_register[6][11] ), .ZN(n1803) );
  INV_X1 U2381 ( .A(\bank_register[18][11] ), .ZN(n1807) );
  INV_X1 U2382 ( .A(\bank_register[7][11] ), .ZN(n1793) );
  INV_X1 U2383 ( .A(\bank_register[19][11] ), .ZN(n1797) );
  INV_X1 U2384 ( .A(\bank_register[6][12] ), .ZN(n1766) );
  INV_X1 U2385 ( .A(\bank_register[18][12] ), .ZN(n1770) );
  INV_X1 U2386 ( .A(\bank_register[7][12] ), .ZN(n1756) );
  INV_X1 U2387 ( .A(\bank_register[19][12] ), .ZN(n1760) );
  INV_X1 U2388 ( .A(\bank_register[6][13] ), .ZN(n1729) );
  INV_X1 U2389 ( .A(\bank_register[18][13] ), .ZN(n1733) );
  INV_X1 U2390 ( .A(\bank_register[7][13] ), .ZN(n1719) );
  INV_X1 U2391 ( .A(\bank_register[19][13] ), .ZN(n1723) );
  INV_X1 U2392 ( .A(\bank_register[6][14] ), .ZN(n1692) );
  INV_X1 U2393 ( .A(\bank_register[18][14] ), .ZN(n1696) );
  INV_X1 U2394 ( .A(\bank_register[7][14] ), .ZN(n1682) );
  INV_X1 U2395 ( .A(\bank_register[19][14] ), .ZN(n1686) );
  INV_X1 U2396 ( .A(\bank_register[6][15] ), .ZN(n1655) );
  INV_X1 U2397 ( .A(\bank_register[18][15] ), .ZN(n1659) );
  INV_X1 U2398 ( .A(\bank_register[7][15] ), .ZN(n1645) );
  INV_X1 U2399 ( .A(\bank_register[19][15] ), .ZN(n1649) );
  INV_X1 U2400 ( .A(\bank_register[6][16] ), .ZN(n1618) );
  INV_X1 U2401 ( .A(\bank_register[18][16] ), .ZN(n1622) );
  INV_X1 U2402 ( .A(\bank_register[7][16] ), .ZN(n1608) );
  INV_X1 U2403 ( .A(\bank_register[19][16] ), .ZN(n1612) );
  INV_X1 U2404 ( .A(\bank_register[6][17] ), .ZN(n1581) );
  INV_X1 U2405 ( .A(\bank_register[18][17] ), .ZN(n1585) );
  INV_X1 U2406 ( .A(\bank_register[7][17] ), .ZN(n1571) );
  INV_X1 U2407 ( .A(\bank_register[19][17] ), .ZN(n1575) );
  INV_X1 U2408 ( .A(\bank_register[6][18] ), .ZN(n1544) );
  INV_X1 U2409 ( .A(\bank_register[18][18] ), .ZN(n1548) );
  INV_X1 U2410 ( .A(\bank_register[7][18] ), .ZN(n1534) );
  INV_X1 U2411 ( .A(\bank_register[19][18] ), .ZN(n1538) );
  INV_X1 U2412 ( .A(\bank_register[6][19] ), .ZN(n1507) );
  INV_X1 U2413 ( .A(\bank_register[18][19] ), .ZN(n1511) );
  INV_X1 U2414 ( .A(\bank_register[7][19] ), .ZN(n1497) );
  INV_X1 U2415 ( .A(\bank_register[19][19] ), .ZN(n1501) );
  INV_X1 U2416 ( .A(\bank_register[6][20] ), .ZN(n1433) );
  INV_X1 U2417 ( .A(\bank_register[18][20] ), .ZN(n1437) );
  INV_X1 U2418 ( .A(\bank_register[7][20] ), .ZN(n1423) );
  INV_X1 U2419 ( .A(\bank_register[19][20] ), .ZN(n1427) );
  INV_X1 U2420 ( .A(\bank_register[6][21] ), .ZN(n1396) );
  INV_X1 U2421 ( .A(\bank_register[18][21] ), .ZN(n1400) );
  INV_X1 U2422 ( .A(\bank_register[7][21] ), .ZN(n1386) );
  INV_X1 U2423 ( .A(\bank_register[19][21] ), .ZN(n1390) );
  INV_X1 U2424 ( .A(\bank_register[6][22] ), .ZN(n1359) );
  INV_X1 U2425 ( .A(\bank_register[18][22] ), .ZN(n1363) );
  INV_X1 U2426 ( .A(\bank_register[7][22] ), .ZN(n1349) );
  INV_X1 U2427 ( .A(\bank_register[19][22] ), .ZN(n1353) );
  INV_X1 U2428 ( .A(\bank_register[6][23] ), .ZN(n1322) );
  INV_X1 U2429 ( .A(\bank_register[18][23] ), .ZN(n1326) );
  INV_X1 U2430 ( .A(\bank_register[7][23] ), .ZN(n1312) );
  INV_X1 U2431 ( .A(\bank_register[19][23] ), .ZN(n1316) );
  INV_X1 U2432 ( .A(\bank_register[6][24] ), .ZN(n1285) );
  INV_X1 U2433 ( .A(\bank_register[18][24] ), .ZN(n1289) );
  INV_X1 U2434 ( .A(\bank_register[7][24] ), .ZN(n1275) );
  INV_X1 U2435 ( .A(\bank_register[19][24] ), .ZN(n1279) );
  INV_X1 U2436 ( .A(\bank_register[6][25] ), .ZN(n1248) );
  INV_X1 U2437 ( .A(\bank_register[18][25] ), .ZN(n1252) );
  INV_X1 U2438 ( .A(\bank_register[7][25] ), .ZN(n1238) );
  INV_X1 U2439 ( .A(\bank_register[19][25] ), .ZN(n1242) );
  INV_X1 U2440 ( .A(\bank_register[6][26] ), .ZN(n1211) );
  INV_X1 U2441 ( .A(\bank_register[18][26] ), .ZN(n1215) );
  INV_X1 U2442 ( .A(\bank_register[7][26] ), .ZN(n1201) );
  INV_X1 U2443 ( .A(\bank_register[19][26] ), .ZN(n1205) );
  INV_X1 U2444 ( .A(\bank_register[6][27] ), .ZN(n1174) );
  INV_X1 U2445 ( .A(\bank_register[18][27] ), .ZN(n1178) );
  INV_X1 U2446 ( .A(\bank_register[7][27] ), .ZN(n1164) );
  INV_X1 U2447 ( .A(\bank_register[19][27] ), .ZN(n1168) );
  INV_X1 U2448 ( .A(\bank_register[6][28] ), .ZN(n1137) );
  INV_X1 U2449 ( .A(\bank_register[18][28] ), .ZN(n1141) );
  INV_X1 U2450 ( .A(\bank_register[7][28] ), .ZN(n1127) );
  INV_X1 U2451 ( .A(\bank_register[19][28] ), .ZN(n1131) );
  INV_X1 U2452 ( .A(\bank_register[6][29] ), .ZN(n1100) );
  INV_X1 U2453 ( .A(\bank_register[18][29] ), .ZN(n1104) );
  INV_X1 U2454 ( .A(\bank_register[7][29] ), .ZN(n1090) );
  INV_X1 U2455 ( .A(\bank_register[19][29] ), .ZN(n1094) );
  INV_X1 U2456 ( .A(\bank_register[6][30] ), .ZN(n1026) );
  INV_X1 U2457 ( .A(\bank_register[18][30] ), .ZN(n1030) );
  INV_X1 U2458 ( .A(\bank_register[7][30] ), .ZN(n1016) );
  INV_X1 U2459 ( .A(\bank_register[19][30] ), .ZN(n1020) );
  INV_X1 U2460 ( .A(\bank_register[6][31] ), .ZN(n989) );
  INV_X1 U2461 ( .A(\bank_register[18][31] ), .ZN(n993) );
  INV_X1 U2462 ( .A(\bank_register[7][31] ), .ZN(n979) );
  INV_X1 U2463 ( .A(\bank_register[19][31] ), .ZN(n983) );
  AND2_X1 U2464 ( .A1(write_data[24]), .A2(n3046), .ZN(n2173) );
  AND2_X1 U2465 ( .A1(write_data[25]), .A2(n3046), .ZN(n2170) );
  AND2_X1 U2466 ( .A1(write_data[26]), .A2(n3046), .ZN(n2167) );
  AND2_X1 U2467 ( .A1(write_data[27]), .A2(n3046), .ZN(n2164) );
  AND2_X1 U2468 ( .A1(write_data[28]), .A2(n3046), .ZN(n2161) );
  AND2_X1 U2469 ( .A1(write_data[29]), .A2(n3046), .ZN(n2158) );
  AND2_X1 U2470 ( .A1(write_data[30]), .A2(n3046), .ZN(n2155) );
  AND2_X1 U2471 ( .A1(write_data[31]), .A2(n3046), .ZN(n2152) );
  AND2_X1 U2472 ( .A1(write_data[6]), .A2(n3047), .ZN(n2227) );
  AND2_X1 U2473 ( .A1(write_data[7]), .A2(n3047), .ZN(n2224) );
  AND2_X1 U2474 ( .A1(write_data[8]), .A2(n3047), .ZN(n2221) );
  AND2_X1 U2475 ( .A1(write_data[9]), .A2(n3047), .ZN(n2218) );
  AND2_X1 U2476 ( .A1(write_data[10]), .A2(n3047), .ZN(n2215) );
  AND2_X1 U2477 ( .A1(write_data[11]), .A2(n3047), .ZN(n2212) );
  AND2_X1 U2478 ( .A1(write_data[12]), .A2(n3047), .ZN(n2209) );
  AND2_X1 U2479 ( .A1(write_data[13]), .A2(n3047), .ZN(n2206) );
  AND2_X1 U2480 ( .A1(write_data[14]), .A2(n3047), .ZN(n2203) );
  AND2_X1 U2481 ( .A1(write_data[15]), .A2(n3047), .ZN(n2200) );
  AND2_X1 U2482 ( .A1(write_data[16]), .A2(n3047), .ZN(n2197) );
  AND2_X1 U2483 ( .A1(write_data[17]), .A2(n3047), .ZN(n2194) );
  AND2_X1 U2484 ( .A1(write_data[18]), .A2(n3047), .ZN(n2191) );
  AND2_X1 U2485 ( .A1(write_data[19]), .A2(n3047), .ZN(n2188) );
  AND2_X1 U2486 ( .A1(write_data[20]), .A2(n3047), .ZN(n2185) );
  AND2_X1 U2487 ( .A1(write_data[21]), .A2(n3047), .ZN(n2182) );
  AND2_X1 U2488 ( .A1(write_data[22]), .A2(n3047), .ZN(n2179) );
  AND2_X1 U2489 ( .A1(write_data[23]), .A2(n3047), .ZN(n2176) );
  AND2_X1 U2490 ( .A1(write_data[0]), .A2(n3048), .ZN(n2245) );
  AND2_X1 U2491 ( .A1(write_data[1]), .A2(n3048), .ZN(n2242) );
  AND2_X1 U2492 ( .A1(write_data[2]), .A2(n3048), .ZN(n2239) );
  AND2_X1 U2493 ( .A1(write_data[3]), .A2(n3048), .ZN(n2236) );
  AND2_X1 U2494 ( .A1(write_data[4]), .A2(n3048), .ZN(n2233) );
  AND2_X1 U2495 ( .A1(write_data[5]), .A2(n3048), .ZN(n2230) );
  INV_X1 U2496 ( .A(\bank_register[20][0] ), .ZN(n2777) );
  INV_X1 U2497 ( .A(\bank_register[24][0] ), .ZN(n2790) );
  INV_X1 U2498 ( .A(\bank_register[20][1] ), .ZN(n2499) );
  INV_X1 U2499 ( .A(\bank_register[24][1] ), .ZN(n2507) );
  INV_X1 U2500 ( .A(\bank_register[20][2] ), .ZN(n2166) );
  INV_X1 U2501 ( .A(\bank_register[24][2] ), .ZN(n2178) );
  INV_X1 U2502 ( .A(\bank_register[20][3] ), .ZN(n2086) );
  INV_X1 U2503 ( .A(\bank_register[24][3] ), .ZN(n2094) );
  INV_X1 U2504 ( .A(\bank_register[20][4] ), .ZN(n2061) );
  INV_X1 U2505 ( .A(\bank_register[24][4] ), .ZN(n2069) );
  INV_X1 U2506 ( .A(\bank_register[20][5] ), .ZN(n2036) );
  INV_X1 U2507 ( .A(\bank_register[24][5] ), .ZN(n2044) );
  INV_X1 U2508 ( .A(\bank_register[20][6] ), .ZN(n2011) );
  INV_X1 U2509 ( .A(\bank_register[24][6] ), .ZN(n2019) );
  INV_X1 U2510 ( .A(\bank_register[20][7] ), .ZN(n1986) );
  INV_X1 U2511 ( .A(\bank_register[24][7] ), .ZN(n1994) );
  INV_X1 U2512 ( .A(\bank_register[20][8] ), .ZN(n1961) );
  INV_X1 U2513 ( .A(\bank_register[24][8] ), .ZN(n1969) );
  INV_X1 U2514 ( .A(\bank_register[20][9] ), .ZN(n1929) );
  INV_X1 U2515 ( .A(\bank_register[24][9] ), .ZN(n1940) );
  INV_X1 U2516 ( .A(\bank_register[20][10] ), .ZN(n2749) );
  INV_X1 U2517 ( .A(\bank_register[24][10] ), .ZN(n2757) );
  INV_X1 U2518 ( .A(\bank_register[20][11] ), .ZN(n2724) );
  INV_X1 U2519 ( .A(\bank_register[24][11] ), .ZN(n2732) );
  INV_X1 U2520 ( .A(\bank_register[20][12] ), .ZN(n2699) );
  INV_X1 U2521 ( .A(\bank_register[24][12] ), .ZN(n2707) );
  INV_X1 U2522 ( .A(\bank_register[20][13] ), .ZN(n2674) );
  INV_X1 U2523 ( .A(\bank_register[24][13] ), .ZN(n2682) );
  INV_X1 U2524 ( .A(\bank_register[20][14] ), .ZN(n2649) );
  INV_X1 U2525 ( .A(\bank_register[24][14] ), .ZN(n2657) );
  INV_X1 U2526 ( .A(\bank_register[20][15] ), .ZN(n2624) );
  INV_X1 U2527 ( .A(\bank_register[24][15] ), .ZN(n2632) );
  INV_X1 U2528 ( .A(\bank_register[20][16] ), .ZN(n2599) );
  INV_X1 U2529 ( .A(\bank_register[24][16] ), .ZN(n2607) );
  INV_X1 U2530 ( .A(\bank_register[20][17] ), .ZN(n2574) );
  INV_X1 U2531 ( .A(\bank_register[24][17] ), .ZN(n2582) );
  INV_X1 U2532 ( .A(\bank_register[20][18] ), .ZN(n2549) );
  INV_X1 U2533 ( .A(\bank_register[24][18] ), .ZN(n2557) );
  INV_X1 U2534 ( .A(\bank_register[20][19] ), .ZN(n2524) );
  INV_X1 U2535 ( .A(\bank_register[24][19] ), .ZN(n2532) );
  INV_X1 U2536 ( .A(\bank_register[20][20] ), .ZN(n2474) );
  INV_X1 U2537 ( .A(\bank_register[24][20] ), .ZN(n2482) );
  INV_X1 U2538 ( .A(\bank_register[20][21] ), .ZN(n2449) );
  INV_X1 U2539 ( .A(\bank_register[24][21] ), .ZN(n2457) );
  INV_X1 U2540 ( .A(\bank_register[20][22] ), .ZN(n2424) );
  INV_X1 U2541 ( .A(\bank_register[24][22] ), .ZN(n2432) );
  INV_X1 U2542 ( .A(\bank_register[20][23] ), .ZN(n2399) );
  INV_X1 U2543 ( .A(\bank_register[24][23] ), .ZN(n2407) );
  INV_X1 U2544 ( .A(\bank_register[20][24] ), .ZN(n2374) );
  INV_X1 U2545 ( .A(\bank_register[24][24] ), .ZN(n2382) );
  INV_X1 U2546 ( .A(\bank_register[20][25] ), .ZN(n2342) );
  INV_X1 U2547 ( .A(\bank_register[24][25] ), .ZN(n2352) );
  INV_X1 U2548 ( .A(\bank_register[20][26] ), .ZN(n2308) );
  INV_X1 U2549 ( .A(\bank_register[24][26] ), .ZN(n2319) );
  INV_X1 U2550 ( .A(\bank_register[20][27] ), .ZN(n2275) );
  INV_X1 U2551 ( .A(\bank_register[24][27] ), .ZN(n2286) );
  INV_X1 U2552 ( .A(\bank_register[20][28] ), .ZN(n2241) );
  INV_X1 U2553 ( .A(\bank_register[24][28] ), .ZN(n2252) );
  INV_X1 U2554 ( .A(\bank_register[20][29] ), .ZN(n2204) );
  INV_X1 U2555 ( .A(\bank_register[24][29] ), .ZN(n2216) );
  INV_X1 U2556 ( .A(\bank_register[20][30] ), .ZN(n2136) );
  INV_X1 U2557 ( .A(\bank_register[24][30] ), .ZN(n2144) );
  INV_X1 U2558 ( .A(\bank_register[20][31] ), .ZN(n2111) );
  INV_X1 U2559 ( .A(\bank_register[24][31] ), .ZN(n2119) );
  INV_X1 U2560 ( .A(\bank_register[28][0] ), .ZN(n2778) );
  INV_X1 U2561 ( .A(\bank_register[28][1] ), .ZN(n2500) );
  INV_X1 U2562 ( .A(\bank_register[28][2] ), .ZN(n2168) );
  INV_X1 U2563 ( .A(\bank_register[28][3] ), .ZN(n2087) );
  INV_X1 U2564 ( .A(\bank_register[28][4] ), .ZN(n2062) );
  INV_X1 U2565 ( .A(\bank_register[28][5] ), .ZN(n2037) );
  INV_X1 U2566 ( .A(\bank_register[28][6] ), .ZN(n2012) );
  INV_X1 U2567 ( .A(\bank_register[28][7] ), .ZN(n1987) );
  INV_X1 U2568 ( .A(\bank_register[28][8] ), .ZN(n1962) );
  INV_X1 U2569 ( .A(\bank_register[28][9] ), .ZN(n1931) );
  INV_X1 U2570 ( .A(\bank_register[28][10] ), .ZN(n2750) );
  INV_X1 U2571 ( .A(\bank_register[28][11] ), .ZN(n2725) );
  INV_X1 U2572 ( .A(\bank_register[28][12] ), .ZN(n2700) );
  INV_X1 U2573 ( .A(\bank_register[28][13] ), .ZN(n2675) );
  INV_X1 U2574 ( .A(\bank_register[28][14] ), .ZN(n2650) );
  INV_X1 U2575 ( .A(\bank_register[28][15] ), .ZN(n2625) );
  INV_X1 U2576 ( .A(\bank_register[28][16] ), .ZN(n2600) );
  INV_X1 U2577 ( .A(\bank_register[28][17] ), .ZN(n2575) );
  INV_X1 U2578 ( .A(\bank_register[28][18] ), .ZN(n2550) );
  INV_X1 U2579 ( .A(\bank_register[28][19] ), .ZN(n2525) );
  INV_X1 U2580 ( .A(\bank_register[28][20] ), .ZN(n2475) );
  INV_X1 U2581 ( .A(\bank_register[28][21] ), .ZN(n2450) );
  INV_X1 U2582 ( .A(\bank_register[28][22] ), .ZN(n2425) );
  INV_X1 U2583 ( .A(\bank_register[28][23] ), .ZN(n2400) );
  INV_X1 U2584 ( .A(\bank_register[28][24] ), .ZN(n2375) );
  INV_X1 U2585 ( .A(\bank_register[28][25] ), .ZN(n2343) );
  INV_X1 U2586 ( .A(\bank_register[28][26] ), .ZN(n2310) );
  INV_X1 U2587 ( .A(\bank_register[28][27] ), .ZN(n2276) );
  INV_X1 U2588 ( .A(\bank_register[28][28] ), .ZN(n2243) );
  INV_X1 U2589 ( .A(\bank_register[28][29] ), .ZN(n2205) );
  INV_X1 U2590 ( .A(\bank_register[28][30] ), .ZN(n2137) );
  INV_X1 U2591 ( .A(\bank_register[28][31] ), .ZN(n2112) );
  INV_X1 U2592 ( .A(write_address[4]), .ZN(n675) );
  INV_X1 U2593 ( .A(write_address[3]), .ZN(n673) );
  INV_X1 U2594 ( .A(N4144), .ZN(n664) );
  CLKBUF_X1 U2595 ( .A(n1920), .Z(n2826) );
  CLKBUF_X1 U2596 ( .A(n1920), .Z(n2827) );
  CLKBUF_X1 U2597 ( .A(n1920), .Z(n2828) );
  CLKBUF_X1 U2598 ( .A(n1919), .Z(n2837) );
  CLKBUF_X1 U2599 ( .A(n1919), .Z(n2838) );
  CLKBUF_X1 U2600 ( .A(n1919), .Z(n2839) );
  CLKBUF_X1 U2601 ( .A(n1917), .Z(n2848) );
  CLKBUF_X1 U2602 ( .A(n1917), .Z(n2849) );
  CLKBUF_X1 U2603 ( .A(n1917), .Z(n2850) );
  CLKBUF_X1 U2604 ( .A(n1916), .Z(n2859) );
  CLKBUF_X1 U2605 ( .A(n1916), .Z(n2860) );
  CLKBUF_X1 U2606 ( .A(n1916), .Z(n2861) );
  CLKBUF_X1 U2607 ( .A(n1915), .Z(n2870) );
  CLKBUF_X1 U2608 ( .A(n1915), .Z(n2871) );
  CLKBUF_X1 U2609 ( .A(n1915), .Z(n2872) );
  CLKBUF_X1 U2610 ( .A(n1914), .Z(n2881) );
  CLKBUF_X1 U2611 ( .A(n1914), .Z(n2882) );
  CLKBUF_X1 U2612 ( .A(n1914), .Z(n2883) );
  CLKBUF_X1 U2613 ( .A(n1912), .Z(n2892) );
  CLKBUF_X1 U2614 ( .A(n1912), .Z(n2893) );
  CLKBUF_X1 U2615 ( .A(n1912), .Z(n2894) );
  CLKBUF_X1 U2616 ( .A(n1911), .Z(n2903) );
  CLKBUF_X1 U2617 ( .A(n1911), .Z(n2904) );
  CLKBUF_X1 U2618 ( .A(n1911), .Z(n2905) );
  CLKBUF_X1 U2619 ( .A(n2905), .Z(n2913) );
  CLKBUF_X1 U2620 ( .A(n714), .Z(n2920) );
  CLKBUF_X1 U2621 ( .A(n714), .Z(n2921) );
  CLKBUF_X1 U2622 ( .A(n714), .Z(n2922) );
  CLKBUF_X1 U2623 ( .A(n712), .Z(n2931) );
  CLKBUF_X1 U2624 ( .A(n712), .Z(n2932) );
  CLKBUF_X1 U2625 ( .A(n712), .Z(n2933) );
  CLKBUF_X1 U2626 ( .A(n710), .Z(n2942) );
  CLKBUF_X1 U2627 ( .A(n710), .Z(n2943) );
  CLKBUF_X1 U2628 ( .A(n710), .Z(n2944) );
  CLKBUF_X1 U2629 ( .A(n2944), .Z(n2952) );
  CLKBUF_X1 U2630 ( .A(n709), .Z(n2953) );
  CLKBUF_X1 U2631 ( .A(n709), .Z(n2954) );
  CLKBUF_X1 U2632 ( .A(n709), .Z(n2955) );
  CLKBUF_X1 U2633 ( .A(n707), .Z(n2964) );
  CLKBUF_X1 U2634 ( .A(n707), .Z(n2965) );
  CLKBUF_X1 U2635 ( .A(n707), .Z(n2966) );
  CLKBUF_X1 U2636 ( .A(n705), .Z(n2975) );
  CLKBUF_X1 U2637 ( .A(n705), .Z(n2976) );
  CLKBUF_X1 U2638 ( .A(n705), .Z(n2977) );
  CLKBUF_X1 U2639 ( .A(n703), .Z(n2986) );
  CLKBUF_X1 U2640 ( .A(n703), .Z(n2987) );
  CLKBUF_X1 U2641 ( .A(n703), .Z(n2988) );
  CLKBUF_X1 U2642 ( .A(n2988), .Z(n2996) );
  CLKBUF_X1 U2643 ( .A(n702), .Z(n2997) );
  CLKBUF_X1 U2644 ( .A(n702), .Z(n2998) );
  CLKBUF_X1 U2645 ( .A(n702), .Z(n2999) );
endmodule


module extender ( immediate, unsigned_value, extended );
  input [15:0] immediate;
  output [31:0] extended;
  input unsigned_value;
  wire   \extended[16] , \immediate[15] , \immediate[14] , \immediate[13] ,
         \immediate[12] , \immediate[11] , \immediate[10] , \immediate[9] ,
         \immediate[8] , \immediate[7] , \immediate[6] , \immediate[5] ,
         \immediate[4] , \immediate[3] , \immediate[2] , \immediate[1] ,
         \immediate[0] , n2;
  assign extended[31] = \extended[16] ;
  assign extended[30] = \extended[16] ;
  assign extended[29] = \extended[16] ;
  assign extended[28] = \extended[16] ;
  assign extended[27] = \extended[16] ;
  assign extended[26] = \extended[16] ;
  assign extended[25] = \extended[16] ;
  assign extended[24] = \extended[16] ;
  assign extended[23] = \extended[16] ;
  assign extended[22] = \extended[16] ;
  assign extended[21] = \extended[16] ;
  assign extended[20] = \extended[16] ;
  assign extended[19] = \extended[16] ;
  assign extended[18] = \extended[16] ;
  assign extended[17] = \extended[16] ;
  assign extended[16] = \extended[16] ;
  assign extended[15] = \immediate[15] ;
  assign \immediate[15]  = immediate[15];
  assign extended[14] = \immediate[14] ;
  assign \immediate[14]  = immediate[14];
  assign extended[13] = \immediate[13] ;
  assign \immediate[13]  = immediate[13];
  assign extended[12] = \immediate[12] ;
  assign \immediate[12]  = immediate[12];
  assign extended[11] = \immediate[11] ;
  assign \immediate[11]  = immediate[11];
  assign extended[10] = \immediate[10] ;
  assign \immediate[10]  = immediate[10];
  assign extended[9] = \immediate[9] ;
  assign \immediate[9]  = immediate[9];
  assign extended[8] = \immediate[8] ;
  assign \immediate[8]  = immediate[8];
  assign extended[7] = \immediate[7] ;
  assign \immediate[7]  = immediate[7];
  assign extended[6] = \immediate[6] ;
  assign \immediate[6]  = immediate[6];
  assign extended[5] = \immediate[5] ;
  assign \immediate[5]  = immediate[5];
  assign extended[4] = \immediate[4] ;
  assign \immediate[4]  = immediate[4];
  assign extended[3] = \immediate[3] ;
  assign \immediate[3]  = immediate[3];
  assign extended[2] = \immediate[2] ;
  assign \immediate[2]  = immediate[2];
  assign extended[1] = \immediate[1] ;
  assign \immediate[1]  = immediate[1];
  assign extended[0] = \immediate[0] ;
  assign \immediate[0]  = immediate[0];

  NOR2_X1 U2 ( .A1(unsigned_value), .A2(n2), .ZN(\extended[16] ) );
  INV_X1 U3 ( .A(\immediate[15] ), .ZN(n2) );
endmodule


module sign_extender ( immediate_jump, extended_jump );
  input [25:0] immediate_jump;
  output [31:0] extended_jump;
  wire   extended_jump_31;
  assign extended_jump[31] = extended_jump_31;
  assign extended_jump[30] = extended_jump_31;
  assign extended_jump[29] = extended_jump_31;
  assign extended_jump[28] = extended_jump_31;
  assign extended_jump[27] = extended_jump_31;
  assign extended_jump[26] = extended_jump_31;
  assign extended_jump[25] = extended_jump_31;
  assign extended_jump_31 = immediate_jump[25];
  assign extended_jump[24] = immediate_jump[24];
  assign extended_jump[23] = immediate_jump[23];
  assign extended_jump[22] = immediate_jump[22];
  assign extended_jump[21] = immediate_jump[21];
  assign extended_jump[20] = immediate_jump[20];
  assign extended_jump[19] = immediate_jump[19];
  assign extended_jump[18] = immediate_jump[18];
  assign extended_jump[17] = immediate_jump[17];
  assign extended_jump[16] = immediate_jump[16];
  assign extended_jump[15] = immediate_jump[15];
  assign extended_jump[14] = immediate_jump[14];
  assign extended_jump[13] = immediate_jump[13];
  assign extended_jump[12] = immediate_jump[12];
  assign extended_jump[11] = immediate_jump[11];
  assign extended_jump[10] = immediate_jump[10];
  assign extended_jump[9] = immediate_jump[9];
  assign extended_jump[8] = immediate_jump[8];
  assign extended_jump[7] = immediate_jump[7];
  assign extended_jump[6] = immediate_jump[6];
  assign extended_jump[5] = immediate_jump[5];
  assign extended_jump[4] = immediate_jump[4];
  assign extended_jump[3] = immediate_jump[3];
  assign extended_jump[2] = immediate_jump[2];
  assign extended_jump[1] = immediate_jump[1];
  assign extended_jump[0] = immediate_jump[0];

endmodule


module mux_stall ( cw_from_cu, mux_op, cw_from_mux );
  input [22:0] cw_from_cu;
  output [22:0] cw_from_mux;
  input mux_op;
  wire   n2;

  AND2_X1 U2 ( .A1(cw_from_cu[7]), .A2(n2), .ZN(cw_from_mux[7]) );
  AND2_X1 U3 ( .A1(cw_from_cu[12]), .A2(n2), .ZN(cw_from_mux[12]) );
  AND2_X1 U4 ( .A1(cw_from_cu[16]), .A2(n2), .ZN(cw_from_mux[16]) );
  AND2_X1 U5 ( .A1(cw_from_cu[18]), .A2(n2), .ZN(cw_from_mux[18]) );
  INV_X1 U6 ( .A(mux_op), .ZN(n2) );
  AND2_X1 U7 ( .A1(cw_from_cu[0]), .A2(n2), .ZN(cw_from_mux[0]) );
  AND2_X1 U8 ( .A1(cw_from_cu[1]), .A2(n2), .ZN(cw_from_mux[1]) );
  AND2_X1 U9 ( .A1(cw_from_cu[5]), .A2(n2), .ZN(cw_from_mux[5]) );
  AND2_X1 U10 ( .A1(cw_from_cu[6]), .A2(n2), .ZN(cw_from_mux[6]) );
  AND2_X1 U11 ( .A1(cw_from_cu[8]), .A2(n2), .ZN(cw_from_mux[8]) );
  AND2_X1 U12 ( .A1(cw_from_cu[9]), .A2(n2), .ZN(cw_from_mux[9]) );
  AND2_X1 U13 ( .A1(cw_from_cu[10]), .A2(n2), .ZN(cw_from_mux[10]) );
  AND2_X1 U14 ( .A1(cw_from_cu[13]), .A2(n2), .ZN(cw_from_mux[13]) );
  AND2_X1 U15 ( .A1(cw_from_cu[17]), .A2(n2), .ZN(cw_from_mux[17]) );
  AND2_X1 U16 ( .A1(cw_from_cu[20]), .A2(n2), .ZN(cw_from_mux[20]) );
  AND2_X1 U17 ( .A1(cw_from_cu[22]), .A2(n2), .ZN(cw_from_mux[22]) );
  AND2_X1 U18 ( .A1(cw_from_cu[21]), .A2(n2), .ZN(cw_from_mux[21]) );
  AND2_X1 U19 ( .A1(cw_from_cu[2]), .A2(n2), .ZN(cw_from_mux[2]) );
  AND2_X1 U20 ( .A1(cw_from_cu[3]), .A2(n2), .ZN(cw_from_mux[3]) );
  AND2_X1 U21 ( .A1(cw_from_cu[4]), .A2(n2), .ZN(cw_from_mux[4]) );
  AND2_X1 U22 ( .A1(cw_from_cu[11]), .A2(n2), .ZN(cw_from_mux[11]) );
  AND2_X1 U23 ( .A1(cw_from_cu[14]), .A2(n2), .ZN(cw_from_mux[14]) );
  AND2_X1 U24 ( .A1(cw_from_cu[15]), .A2(n2), .ZN(cw_from_mux[15]) );
  AND2_X1 U25 ( .A1(cw_from_cu[19]), .A2(n2), .ZN(cw_from_mux[19]) );
endmodule


module hdu ( clk, rst, idex_mem_read, idex_rt, rs, rt, pcwrite, ifidwrite, 
        mux_op );
  input [3:0] idex_mem_read;
  input [4:0] idex_rt;
  input [4:0] rs;
  input [4:0] rt;
  input clk, rst;
  output pcwrite, ifidwrite, mux_op;
  wire   ifidwrite, N7, N8, n6, net41391, n7, n8, n9, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;
  assign pcwrite = ifidwrite;

  DFF_X1 \current_state_reg[0]  ( .D(N7), .CK(clk), .QN(net41391) );
  DFF_X1 \current_state_reg[1]  ( .D(N8), .CK(clk), .Q(n6), .QN(n25) );
  OAI33_X1 U18 ( .A1(n13), .A2(n14), .A3(n15), .B1(n16), .B2(n17), .B3(n18), 
        .ZN(n11) );
  XOR2_X1 U19 ( .A(rt[4]), .B(idex_rt[4]), .Z(n18) );
  XOR2_X1 U20 ( .A(rt[2]), .B(idex_rt[2]), .Z(n17) );
  NAND3_X1 U21 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n16) );
  XOR2_X1 U22 ( .A(rs[4]), .B(idex_rt[4]), .Z(n15) );
  XOR2_X1 U23 ( .A(rs[3]), .B(idex_rt[3]), .Z(n14) );
  NAND3_X1 U24 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n13) );
  INV_X1 U3 ( .A(n7), .ZN(ifidwrite) );
  NOR3_X1 U4 ( .A1(n6), .A2(net41391), .A3(n9), .ZN(mux_op) );
  AOI21_X1 U5 ( .B1(n25), .B2(n9), .A(net41391), .ZN(n7) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(n9) );
  OR4_X1 U7 ( .A1(idex_mem_read[1]), .A2(idex_mem_read[0]), .A3(
        idex_mem_read[3]), .A4(idex_mem_read[2]), .ZN(n12) );
  XNOR2_X1 U8 ( .A(idex_rt[0]), .B(rs[0]), .ZN(n22) );
  XNOR2_X1 U9 ( .A(idex_rt[1]), .B(rs[1]), .ZN(n23) );
  XNOR2_X1 U10 ( .A(idex_rt[2]), .B(rs[2]), .ZN(n24) );
  XNOR2_X1 U11 ( .A(idex_rt[0]), .B(rt[0]), .ZN(n20) );
  XNOR2_X1 U12 ( .A(idex_rt[3]), .B(rt[3]), .ZN(n19) );
  XNOR2_X1 U13 ( .A(idex_rt[1]), .B(rt[1]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(rst), .A2(n7), .ZN(N7) );
  NOR2_X1 U15 ( .A1(rst), .A2(n8), .ZN(N8) );
  INV_X1 U16 ( .A(mux_op), .ZN(n8) );
endmodule


module iram_block ( from_pc, flush, from_iram, to_iram, to_if_id_reg );
  input [31:0] from_pc;
  input [31:0] from_iram;
  output [31:0] to_iram;
  output [31:0] to_if_id_reg;
  input flush;

  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign to_iram[31] = 1'b0;
  assign to_iram[30] = 1'b0;

  mmu_in_iram mmu_in ( .from_pc(from_pc), .to_iram({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, to_iram[29:0]}) );
  mmu_out_iram mmu_out ( .from_iram(from_iram), .flush(flush), .to_if_id_reg(
        to_if_id_reg) );
endmodule


module increment_pc ( from_pc, to_mux_branch );
  input [31:0] from_pc;
  output [31:0] to_mux_branch;


  increment_pc_DW01_add_0 add_33 ( .A(from_pc), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(to_mux_branch) );
endmodule


module pc ( from_mux_jump, pcwrite, clk, rst, to_iram_block );
  input [31:0] from_mux_jump;
  output [31:0] to_iram_block;
  input pcwrite, clk, rst;
  wire   n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n34, n35, n36, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138;

  DFF_X1 \to_iram_block_reg[31]  ( .D(n100), .CK(clk), .Q(to_iram_block[31]), 
        .QN(n37) );
  DFF_X1 \to_iram_block_reg[30]  ( .D(n99), .CK(clk), .Q(to_iram_block[30]), 
        .QN(n38) );
  DFF_X1 \to_iram_block_reg[29]  ( .D(n98), .CK(clk), .Q(to_iram_block[29]), 
        .QN(n39) );
  DFF_X1 \to_iram_block_reg[28]  ( .D(n97), .CK(clk), .Q(to_iram_block[28]), 
        .QN(n40) );
  DFF_X1 \to_iram_block_reg[27]  ( .D(n96), .CK(clk), .Q(to_iram_block[27]), 
        .QN(n41) );
  DFF_X1 \to_iram_block_reg[26]  ( .D(n95), .CK(clk), .Q(to_iram_block[26]), 
        .QN(n42) );
  DFF_X1 \to_iram_block_reg[25]  ( .D(n94), .CK(clk), .Q(to_iram_block[25]), 
        .QN(n43) );
  DFF_X1 \to_iram_block_reg[24]  ( .D(n93), .CK(clk), .Q(to_iram_block[24]), 
        .QN(n44) );
  DFF_X1 \to_iram_block_reg[23]  ( .D(n92), .CK(clk), .Q(to_iram_block[23]), 
        .QN(n45) );
  DFF_X1 \to_iram_block_reg[22]  ( .D(n91), .CK(clk), .Q(to_iram_block[22]), 
        .QN(n46) );
  DFF_X1 \to_iram_block_reg[21]  ( .D(n90), .CK(clk), .Q(to_iram_block[21]), 
        .QN(n47) );
  DFF_X1 \to_iram_block_reg[20]  ( .D(n89), .CK(clk), .Q(to_iram_block[20]), 
        .QN(n48) );
  DFF_X1 \to_iram_block_reg[19]  ( .D(n88), .CK(clk), .Q(to_iram_block[19]), 
        .QN(n49) );
  DFF_X1 \to_iram_block_reg[18]  ( .D(n87), .CK(clk), .Q(to_iram_block[18]), 
        .QN(n50) );
  DFF_X1 \to_iram_block_reg[17]  ( .D(n86), .CK(clk), .Q(to_iram_block[17]), 
        .QN(n51) );
  DFF_X1 \to_iram_block_reg[16]  ( .D(n85), .CK(clk), .Q(to_iram_block[16]), 
        .QN(n52) );
  DFF_X1 \to_iram_block_reg[15]  ( .D(n84), .CK(clk), .Q(to_iram_block[15]), 
        .QN(n53) );
  DFF_X1 \to_iram_block_reg[14]  ( .D(n83), .CK(clk), .Q(to_iram_block[14]), 
        .QN(n54) );
  DFF_X1 \to_iram_block_reg[13]  ( .D(n82), .CK(clk), .Q(to_iram_block[13]), 
        .QN(n55) );
  DFF_X1 \to_iram_block_reg[12]  ( .D(n81), .CK(clk), .Q(to_iram_block[12]), 
        .QN(n56) );
  DFF_X1 \to_iram_block_reg[11]  ( .D(n80), .CK(clk), .Q(to_iram_block[11]), 
        .QN(n57) );
  DFF_X1 \to_iram_block_reg[10]  ( .D(n79), .CK(clk), .Q(to_iram_block[10]), 
        .QN(n58) );
  DFF_X1 \to_iram_block_reg[9]  ( .D(n78), .CK(clk), .Q(to_iram_block[9]), 
        .QN(n59) );
  DFF_X1 \to_iram_block_reg[8]  ( .D(n77), .CK(clk), .Q(to_iram_block[8]), 
        .QN(n60) );
  DFF_X1 \to_iram_block_reg[7]  ( .D(n76), .CK(clk), .Q(to_iram_block[7]), 
        .QN(n61) );
  DFF_X1 \to_iram_block_reg[6]  ( .D(n75), .CK(clk), .Q(to_iram_block[6]), 
        .QN(n62) );
  DFF_X1 \to_iram_block_reg[5]  ( .D(n74), .CK(clk), .Q(to_iram_block[5]), 
        .QN(n63) );
  DFF_X1 \to_iram_block_reg[4]  ( .D(n73), .CK(clk), .Q(to_iram_block[4]), 
        .QN(n64) );
  DFF_X1 \to_iram_block_reg[3]  ( .D(n72), .CK(clk), .Q(to_iram_block[3]), 
        .QN(n65) );
  DFF_X1 \to_iram_block_reg[2]  ( .D(n71), .CK(clk), .Q(to_iram_block[2]), 
        .QN(n66) );
  DFF_X1 \to_iram_block_reg[1]  ( .D(n70), .CK(clk), .Q(to_iram_block[1]), 
        .QN(n67) );
  DFF_X1 \to_iram_block_reg[0]  ( .D(n69), .CK(clk), .Q(to_iram_block[0]), 
        .QN(n68) );
  BUF_X1 U3 ( .A(n34), .Z(n136) );
  BUF_X1 U4 ( .A(n34), .Z(n137) );
  BUF_X1 U5 ( .A(n35), .Z(n134) );
  BUF_X1 U6 ( .A(n35), .Z(n133) );
  BUF_X1 U7 ( .A(n35), .Z(n135) );
  BUF_X1 U8 ( .A(n34), .Z(n138) );
  OAI22_X1 U9 ( .A1(n137), .A2(n45), .B1(n135), .B2(n107), .ZN(n92) );
  INV_X1 U10 ( .A(from_mux_jump[23]), .ZN(n107) );
  OAI22_X1 U11 ( .A1(n138), .A2(n44), .B1(n135), .B2(n106), .ZN(n93) );
  INV_X1 U12 ( .A(from_mux_jump[24]), .ZN(n106) );
  OAI22_X1 U13 ( .A1(n138), .A2(n41), .B1(n135), .B2(n103), .ZN(n96) );
  INV_X1 U14 ( .A(from_mux_jump[27]), .ZN(n103) );
  OAI22_X1 U15 ( .A1(n138), .A2(n40), .B1(n135), .B2(n102), .ZN(n97) );
  INV_X1 U16 ( .A(from_mux_jump[28]), .ZN(n102) );
  OAI22_X1 U17 ( .A1(n137), .A2(n53), .B1(n134), .B2(n115), .ZN(n84) );
  INV_X1 U18 ( .A(from_mux_jump[15]), .ZN(n115) );
  OAI22_X1 U19 ( .A1(n137), .A2(n52), .B1(n134), .B2(n114), .ZN(n85) );
  INV_X1 U20 ( .A(from_mux_jump[16]), .ZN(n114) );
  OAI22_X1 U21 ( .A1(n137), .A2(n49), .B1(n134), .B2(n111), .ZN(n88) );
  INV_X1 U22 ( .A(from_mux_jump[19]), .ZN(n111) );
  OAI22_X1 U23 ( .A1(n136), .A2(n37), .B1(n133), .B2(n131), .ZN(n100) );
  INV_X1 U24 ( .A(from_mux_jump[31]), .ZN(n131) );
  OAI22_X1 U25 ( .A1(n137), .A2(n54), .B1(n134), .B2(n116), .ZN(n83) );
  INV_X1 U26 ( .A(from_mux_jump[14]), .ZN(n116) );
  OAI22_X1 U27 ( .A1(n137), .A2(n51), .B1(n134), .B2(n113), .ZN(n86) );
  INV_X1 U28 ( .A(from_mux_jump[17]), .ZN(n113) );
  OAI22_X1 U29 ( .A1(n137), .A2(n50), .B1(n134), .B2(n112), .ZN(n87) );
  INV_X1 U30 ( .A(from_mux_jump[18]), .ZN(n112) );
  OAI22_X1 U31 ( .A1(n137), .A2(n48), .B1(n134), .B2(n110), .ZN(n89) );
  INV_X1 U32 ( .A(from_mux_jump[20]), .ZN(n110) );
  OAI22_X1 U33 ( .A1(n137), .A2(n47), .B1(n134), .B2(n109), .ZN(n90) );
  INV_X1 U34 ( .A(from_mux_jump[21]), .ZN(n109) );
  OAI22_X1 U35 ( .A1(n137), .A2(n46), .B1(n134), .B2(n108), .ZN(n91) );
  INV_X1 U36 ( .A(from_mux_jump[22]), .ZN(n108) );
  OAI22_X1 U37 ( .A1(n138), .A2(n43), .B1(n135), .B2(n105), .ZN(n94) );
  INV_X1 U38 ( .A(from_mux_jump[25]), .ZN(n105) );
  OAI22_X1 U39 ( .A1(n138), .A2(n42), .B1(n135), .B2(n104), .ZN(n95) );
  INV_X1 U40 ( .A(from_mux_jump[26]), .ZN(n104) );
  OAI22_X1 U41 ( .A1(n138), .A2(n39), .B1(n135), .B2(n101), .ZN(n98) );
  INV_X1 U42 ( .A(from_mux_jump[29]), .ZN(n101) );
  OAI22_X1 U43 ( .A1(n138), .A2(n38), .B1(n135), .B2(n36), .ZN(n99) );
  INV_X1 U44 ( .A(from_mux_jump[30]), .ZN(n36) );
  OAI22_X1 U45 ( .A1(n136), .A2(n68), .B1(n133), .B2(n130), .ZN(n69) );
  INV_X1 U46 ( .A(from_mux_jump[0]), .ZN(n130) );
  OAI22_X1 U47 ( .A1(n136), .A2(n67), .B1(n133), .B2(n129), .ZN(n70) );
  INV_X1 U48 ( .A(from_mux_jump[1]), .ZN(n129) );
  OAI22_X1 U49 ( .A1(n136), .A2(n66), .B1(n133), .B2(n128), .ZN(n71) );
  INV_X1 U50 ( .A(from_mux_jump[2]), .ZN(n128) );
  OAI22_X1 U51 ( .A1(n136), .A2(n65), .B1(n133), .B2(n127), .ZN(n72) );
  INV_X1 U52 ( .A(from_mux_jump[3]), .ZN(n127) );
  OAI22_X1 U53 ( .A1(n136), .A2(n64), .B1(n133), .B2(n126), .ZN(n73) );
  INV_X1 U54 ( .A(from_mux_jump[4]), .ZN(n126) );
  OAI22_X1 U55 ( .A1(n136), .A2(n63), .B1(n133), .B2(n125), .ZN(n74) );
  INV_X1 U56 ( .A(from_mux_jump[5]), .ZN(n125) );
  OAI22_X1 U57 ( .A1(n136), .A2(n62), .B1(n133), .B2(n124), .ZN(n75) );
  INV_X1 U58 ( .A(from_mux_jump[6]), .ZN(n124) );
  OAI22_X1 U59 ( .A1(n136), .A2(n61), .B1(n133), .B2(n123), .ZN(n76) );
  INV_X1 U60 ( .A(from_mux_jump[7]), .ZN(n123) );
  OAI22_X1 U61 ( .A1(n136), .A2(n60), .B1(n133), .B2(n122), .ZN(n77) );
  INV_X1 U62 ( .A(from_mux_jump[8]), .ZN(n122) );
  OAI22_X1 U63 ( .A1(n136), .A2(n59), .B1(n133), .B2(n121), .ZN(n78) );
  INV_X1 U64 ( .A(from_mux_jump[9]), .ZN(n121) );
  OAI22_X1 U65 ( .A1(n136), .A2(n58), .B1(n133), .B2(n120), .ZN(n79) );
  INV_X1 U66 ( .A(from_mux_jump[10]), .ZN(n120) );
  OAI22_X1 U67 ( .A1(n137), .A2(n57), .B1(n134), .B2(n119), .ZN(n80) );
  INV_X1 U68 ( .A(from_mux_jump[11]), .ZN(n119) );
  OAI22_X1 U69 ( .A1(n137), .A2(n56), .B1(n134), .B2(n118), .ZN(n81) );
  INV_X1 U70 ( .A(from_mux_jump[12]), .ZN(n118) );
  NAND2_X1 U71 ( .A1(n132), .A2(n136), .ZN(n35) );
  INV_X1 U72 ( .A(rst), .ZN(n132) );
  OR2_X1 U73 ( .A1(pcwrite), .A2(rst), .ZN(n34) );
  OAI22_X1 U74 ( .A1(n137), .A2(n55), .B1(n134), .B2(n117), .ZN(n82) );
  INV_X1 U75 ( .A(from_mux_jump[13]), .ZN(n117) );
endmodule


module mux_jump ( jump_address, from_mux_branch, jump, to_pc );
  input [31:0] jump_address;
  input [31:0] from_mux_branch;
  output [31:0] to_pc;
  input jump;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28;

  INV_X1 U1 ( .A(n28), .ZN(n18) );
  INV_X1 U2 ( .A(n28), .ZN(n19) );
  BUF_X1 U3 ( .A(n15), .Z(n20) );
  BUF_X1 U4 ( .A(n17), .Z(n27) );
  BUF_X1 U5 ( .A(n17), .Z(n26) );
  BUF_X1 U6 ( .A(n16), .Z(n25) );
  BUF_X1 U7 ( .A(n16), .Z(n24) );
  BUF_X1 U8 ( .A(n16), .Z(n23) );
  BUF_X1 U9 ( .A(n15), .Z(n22) );
  BUF_X1 U10 ( .A(n15), .Z(n21) );
  BUF_X1 U11 ( .A(n17), .Z(n28) );
  INV_X1 U12 ( .A(n51), .ZN(to_pc[23]) );
  AOI22_X1 U13 ( .A1(from_mux_branch[23]), .A2(n19), .B1(jump_address[23]), 
        .B2(n24), .ZN(n51) );
  INV_X1 U14 ( .A(n50), .ZN(to_pc[24]) );
  AOI22_X1 U15 ( .A1(from_mux_branch[24]), .A2(n19), .B1(jump_address[24]), 
        .B2(n23), .ZN(n50) );
  INV_X1 U16 ( .A(n47), .ZN(to_pc[27]) );
  AOI22_X1 U17 ( .A1(from_mux_branch[27]), .A2(n19), .B1(jump_address[27]), 
        .B2(n23), .ZN(n47) );
  INV_X1 U18 ( .A(n46), .ZN(to_pc[28]) );
  AOI22_X1 U19 ( .A1(from_mux_branch[28]), .A2(n19), .B1(jump_address[28]), 
        .B2(n22), .ZN(n46) );
  INV_X1 U20 ( .A(n60), .ZN(to_pc[15]) );
  AOI22_X1 U21 ( .A1(from_mux_branch[15]), .A2(n18), .B1(jump_address[15]), 
        .B2(n26), .ZN(n60) );
  INV_X1 U22 ( .A(n59), .ZN(to_pc[16]) );
  AOI22_X1 U23 ( .A1(from_mux_branch[16]), .A2(n18), .B1(jump_address[16]), 
        .B2(n26), .ZN(n59) );
  INV_X1 U24 ( .A(n56), .ZN(to_pc[19]) );
  AOI22_X1 U25 ( .A1(from_mux_branch[19]), .A2(n18), .B1(jump_address[19]), 
        .B2(n25), .ZN(n56) );
  INV_X1 U26 ( .A(n42), .ZN(to_pc[31]) );
  AOI22_X1 U27 ( .A1(from_mux_branch[31]), .A2(n18), .B1(jump_address[31]), 
        .B2(n21), .ZN(n42) );
  INV_X1 U28 ( .A(n61), .ZN(to_pc[14]) );
  AOI22_X1 U29 ( .A1(from_mux_branch[14]), .A2(n18), .B1(jump_address[14]), 
        .B2(n26), .ZN(n61) );
  INV_X1 U30 ( .A(n58), .ZN(to_pc[17]) );
  AOI22_X1 U31 ( .A1(from_mux_branch[17]), .A2(n18), .B1(jump_address[17]), 
        .B2(n25), .ZN(n58) );
  INV_X1 U32 ( .A(n57), .ZN(to_pc[18]) );
  AOI22_X1 U33 ( .A1(from_mux_branch[18]), .A2(n18), .B1(jump_address[18]), 
        .B2(n25), .ZN(n57) );
  INV_X1 U34 ( .A(n54), .ZN(to_pc[20]) );
  AOI22_X1 U35 ( .A1(from_mux_branch[20]), .A2(n19), .B1(jump_address[20]), 
        .B2(n24), .ZN(n54) );
  INV_X1 U36 ( .A(n53), .ZN(to_pc[21]) );
  AOI22_X1 U37 ( .A1(from_mux_branch[21]), .A2(n19), .B1(jump_address[21]), 
        .B2(n24), .ZN(n53) );
  INV_X1 U38 ( .A(n52), .ZN(to_pc[22]) );
  AOI22_X1 U39 ( .A1(from_mux_branch[22]), .A2(n19), .B1(jump_address[22]), 
        .B2(n24), .ZN(n52) );
  INV_X1 U40 ( .A(n49), .ZN(to_pc[25]) );
  AOI22_X1 U41 ( .A1(from_mux_branch[25]), .A2(n19), .B1(jump_address[25]), 
        .B2(n23), .ZN(n49) );
  INV_X1 U42 ( .A(n48), .ZN(to_pc[26]) );
  AOI22_X1 U43 ( .A1(from_mux_branch[26]), .A2(n19), .B1(jump_address[26]), 
        .B2(n23), .ZN(n48) );
  INV_X1 U44 ( .A(n45), .ZN(to_pc[29]) );
  AOI22_X1 U45 ( .A1(from_mux_branch[29]), .A2(n19), .B1(jump_address[29]), 
        .B2(n22), .ZN(n45) );
  INV_X1 U46 ( .A(n43), .ZN(to_pc[30]) );
  AOI22_X1 U47 ( .A1(from_mux_branch[30]), .A2(n19), .B1(jump_address[30]), 
        .B2(n22), .ZN(n43) );
  INV_X1 U48 ( .A(n66), .ZN(to_pc[0]) );
  AOI22_X1 U49 ( .A1(from_mux_branch[0]), .A2(n18), .B1(jump_address[0]), .B2(
        n27), .ZN(n66) );
  INV_X1 U50 ( .A(n55), .ZN(to_pc[1]) );
  AOI22_X1 U51 ( .A1(from_mux_branch[1]), .A2(n18), .B1(jump_address[1]), .B2(
        n25), .ZN(n55) );
  INV_X1 U52 ( .A(n44), .ZN(to_pc[2]) );
  AOI22_X1 U53 ( .A1(from_mux_branch[2]), .A2(n19), .B1(jump_address[2]), .B2(
        n22), .ZN(n44) );
  INV_X1 U54 ( .A(n41), .ZN(to_pc[3]) );
  AOI22_X1 U55 ( .A1(from_mux_branch[3]), .A2(n19), .B1(jump_address[3]), .B2(
        n21), .ZN(n41) );
  INV_X1 U56 ( .A(n40), .ZN(to_pc[4]) );
  AOI22_X1 U57 ( .A1(from_mux_branch[4]), .A2(n18), .B1(jump_address[4]), .B2(
        n21), .ZN(n40) );
  INV_X1 U58 ( .A(n39), .ZN(to_pc[5]) );
  AOI22_X1 U59 ( .A1(from_mux_branch[5]), .A2(n19), .B1(jump_address[5]), .B2(
        n21), .ZN(n39) );
  INV_X1 U60 ( .A(n38), .ZN(to_pc[6]) );
  AOI22_X1 U61 ( .A1(from_mux_branch[6]), .A2(n18), .B1(jump_address[6]), .B2(
        n20), .ZN(n38) );
  INV_X1 U62 ( .A(n37), .ZN(to_pc[7]) );
  AOI22_X1 U63 ( .A1(from_mux_branch[7]), .A2(n19), .B1(jump_address[7]), .B2(
        n20), .ZN(n37) );
  INV_X1 U64 ( .A(n36), .ZN(to_pc[8]) );
  AOI22_X1 U65 ( .A1(from_mux_branch[8]), .A2(n18), .B1(jump_address[8]), .B2(
        n20), .ZN(n36) );
  INV_X1 U66 ( .A(n34), .ZN(to_pc[9]) );
  AOI22_X1 U67 ( .A1(from_mux_branch[9]), .A2(n19), .B1(jump_address[9]), .B2(
        n20), .ZN(n34) );
  INV_X1 U68 ( .A(n65), .ZN(to_pc[10]) );
  AOI22_X1 U69 ( .A1(from_mux_branch[10]), .A2(n18), .B1(jump_address[10]), 
        .B2(n27), .ZN(n65) );
  INV_X1 U70 ( .A(n64), .ZN(to_pc[11]) );
  AOI22_X1 U71 ( .A1(from_mux_branch[11]), .A2(n18), .B1(jump_address[11]), 
        .B2(n27), .ZN(n64) );
  INV_X1 U72 ( .A(n63), .ZN(to_pc[12]) );
  AOI22_X1 U73 ( .A1(from_mux_branch[12]), .A2(n18), .B1(jump_address[12]), 
        .B2(n27), .ZN(n63) );
  BUF_X1 U74 ( .A(jump), .Z(n17) );
  BUF_X1 U75 ( .A(jump), .Z(n16) );
  BUF_X1 U76 ( .A(jump), .Z(n15) );
  INV_X1 U77 ( .A(n62), .ZN(to_pc[13]) );
  AOI22_X1 U78 ( .A1(from_mux_branch[13]), .A2(n18), .B1(jump_address[13]), 
        .B2(n26), .ZN(n62) );
endmodule


module mux_branch ( from_increment_pc, branch_target, pcsrc, to_mux_jump );
  input [31:0] from_increment_pc;
  input [31:0] branch_target;
  output [31:0] to_mux_jump;
  input pcsrc;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22;

  INV_X1 U1 ( .A(n21), .ZN(n12) );
  BUF_X1 U2 ( .A(n22), .Z(n13) );
  BUF_X1 U3 ( .A(n13), .Z(n20) );
  BUF_X1 U4 ( .A(n17), .Z(n19) );
  BUF_X1 U5 ( .A(n22), .Z(n18) );
  BUF_X1 U6 ( .A(n22), .Z(n17) );
  BUF_X1 U7 ( .A(n22), .Z(n16) );
  BUF_X1 U8 ( .A(n22), .Z(n15) );
  BUF_X1 U9 ( .A(n22), .Z(n14) );
  BUF_X1 U10 ( .A(n22), .Z(n21) );
  INV_X1 U11 ( .A(pcsrc), .ZN(n22) );
  INV_X1 U12 ( .A(n61), .ZN(to_mux_jump[14]) );
  AOI22_X1 U13 ( .A1(branch_target[14]), .A2(n12), .B1(from_increment_pc[14]), 
        .B2(n19), .ZN(n61) );
  INV_X1 U14 ( .A(n60), .ZN(to_mux_jump[15]) );
  AOI22_X1 U15 ( .A1(branch_target[15]), .A2(n12), .B1(from_increment_pc[15]), 
        .B2(n19), .ZN(n60) );
  INV_X1 U16 ( .A(n59), .ZN(to_mux_jump[16]) );
  AOI22_X1 U17 ( .A1(branch_target[16]), .A2(n12), .B1(from_increment_pc[16]), 
        .B2(n19), .ZN(n59) );
  INV_X1 U18 ( .A(n58), .ZN(to_mux_jump[17]) );
  AOI22_X1 U19 ( .A1(branch_target[17]), .A2(n12), .B1(from_increment_pc[17]), 
        .B2(n18), .ZN(n58) );
  INV_X1 U20 ( .A(n57), .ZN(to_mux_jump[18]) );
  AOI22_X1 U21 ( .A1(branch_target[18]), .A2(n12), .B1(from_increment_pc[18]), 
        .B2(n18), .ZN(n57) );
  INV_X1 U22 ( .A(n56), .ZN(to_mux_jump[19]) );
  AOI22_X1 U23 ( .A1(branch_target[19]), .A2(n12), .B1(from_increment_pc[19]), 
        .B2(n18), .ZN(n56) );
  INV_X1 U24 ( .A(n54), .ZN(to_mux_jump[20]) );
  AOI22_X1 U25 ( .A1(branch_target[20]), .A2(pcsrc), .B1(from_increment_pc[20]), .B2(n17), .ZN(n54) );
  INV_X1 U26 ( .A(n53), .ZN(to_mux_jump[21]) );
  AOI22_X1 U27 ( .A1(branch_target[21]), .A2(pcsrc), .B1(from_increment_pc[21]), .B2(n17), .ZN(n53) );
  INV_X1 U28 ( .A(n52), .ZN(to_mux_jump[22]) );
  AOI22_X1 U29 ( .A1(branch_target[22]), .A2(n12), .B1(from_increment_pc[22]), 
        .B2(n17), .ZN(n52) );
  INV_X1 U30 ( .A(n51), .ZN(to_mux_jump[23]) );
  AOI22_X1 U31 ( .A1(branch_target[23]), .A2(pcsrc), .B1(from_increment_pc[23]), .B2(n17), .ZN(n51) );
  INV_X1 U32 ( .A(n50), .ZN(to_mux_jump[24]) );
  AOI22_X1 U33 ( .A1(branch_target[24]), .A2(pcsrc), .B1(from_increment_pc[24]), .B2(n16), .ZN(n50) );
  INV_X1 U34 ( .A(n49), .ZN(to_mux_jump[25]) );
  AOI22_X1 U35 ( .A1(branch_target[25]), .A2(pcsrc), .B1(from_increment_pc[25]), .B2(n16), .ZN(n49) );
  INV_X1 U36 ( .A(n48), .ZN(to_mux_jump[26]) );
  AOI22_X1 U37 ( .A1(branch_target[26]), .A2(pcsrc), .B1(from_increment_pc[26]), .B2(n16), .ZN(n48) );
  INV_X1 U38 ( .A(n47), .ZN(to_mux_jump[27]) );
  AOI22_X1 U39 ( .A1(branch_target[27]), .A2(pcsrc), .B1(from_increment_pc[27]), .B2(n16), .ZN(n47) );
  INV_X1 U40 ( .A(n46), .ZN(to_mux_jump[28]) );
  AOI22_X1 U41 ( .A1(branch_target[28]), .A2(pcsrc), .B1(from_increment_pc[28]), .B2(n15), .ZN(n46) );
  INV_X1 U42 ( .A(n45), .ZN(to_mux_jump[29]) );
  AOI22_X1 U43 ( .A1(branch_target[29]), .A2(pcsrc), .B1(from_increment_pc[29]), .B2(n15), .ZN(n45) );
  INV_X1 U44 ( .A(n43), .ZN(to_mux_jump[30]) );
  AOI22_X1 U45 ( .A1(branch_target[30]), .A2(pcsrc), .B1(from_increment_pc[30]), .B2(n15), .ZN(n43) );
  INV_X1 U46 ( .A(n42), .ZN(to_mux_jump[31]) );
  AOI22_X1 U47 ( .A1(branch_target[31]), .A2(pcsrc), .B1(from_increment_pc[31]), .B2(n14), .ZN(n42) );
  INV_X1 U48 ( .A(n34), .ZN(to_mux_jump[9]) );
  AOI22_X1 U49 ( .A1(pcsrc), .A2(branch_target[9]), .B1(from_increment_pc[9]), 
        .B2(n13), .ZN(n34) );
  INV_X1 U50 ( .A(n41), .ZN(to_mux_jump[3]) );
  AOI22_X1 U51 ( .A1(branch_target[3]), .A2(pcsrc), .B1(from_increment_pc[3]), 
        .B2(n14), .ZN(n41) );
  INV_X1 U52 ( .A(n40), .ZN(to_mux_jump[4]) );
  AOI22_X1 U53 ( .A1(branch_target[4]), .A2(pcsrc), .B1(from_increment_pc[4]), 
        .B2(n14), .ZN(n40) );
  INV_X1 U54 ( .A(n39), .ZN(to_mux_jump[5]) );
  AOI22_X1 U55 ( .A1(branch_target[5]), .A2(pcsrc), .B1(from_increment_pc[5]), 
        .B2(n14), .ZN(n39) );
  INV_X1 U56 ( .A(n38), .ZN(to_mux_jump[6]) );
  AOI22_X1 U57 ( .A1(branch_target[6]), .A2(pcsrc), .B1(from_increment_pc[6]), 
        .B2(n13), .ZN(n38) );
  INV_X1 U58 ( .A(n37), .ZN(to_mux_jump[7]) );
  AOI22_X1 U59 ( .A1(branch_target[7]), .A2(n12), .B1(from_increment_pc[7]), 
        .B2(n13), .ZN(n37) );
  INV_X1 U60 ( .A(n36), .ZN(to_mux_jump[8]) );
  AOI22_X1 U61 ( .A1(branch_target[8]), .A2(pcsrc), .B1(from_increment_pc[8]), 
        .B2(n13), .ZN(n36) );
  INV_X1 U62 ( .A(n65), .ZN(to_mux_jump[10]) );
  AOI22_X1 U63 ( .A1(branch_target[10]), .A2(n12), .B1(from_increment_pc[10]), 
        .B2(n20), .ZN(n65) );
  INV_X1 U64 ( .A(n64), .ZN(to_mux_jump[11]) );
  AOI22_X1 U65 ( .A1(branch_target[11]), .A2(n12), .B1(from_increment_pc[11]), 
        .B2(n20), .ZN(n64) );
  INV_X1 U66 ( .A(n63), .ZN(to_mux_jump[12]) );
  AOI22_X1 U67 ( .A1(branch_target[12]), .A2(n12), .B1(from_increment_pc[12]), 
        .B2(n20), .ZN(n63) );
  INV_X1 U68 ( .A(n62), .ZN(to_mux_jump[13]) );
  AOI22_X1 U69 ( .A1(branch_target[13]), .A2(n12), .B1(from_increment_pc[13]), 
        .B2(n19), .ZN(n62) );
  INV_X1 U70 ( .A(n66), .ZN(to_mux_jump[0]) );
  AOI22_X1 U71 ( .A1(branch_target[0]), .A2(n12), .B1(from_increment_pc[0]), 
        .B2(n20), .ZN(n66) );
  INV_X1 U72 ( .A(n55), .ZN(to_mux_jump[1]) );
  AOI22_X1 U73 ( .A1(branch_target[1]), .A2(n12), .B1(from_increment_pc[1]), 
        .B2(n18), .ZN(n55) );
  INV_X1 U74 ( .A(n44), .ZN(to_mux_jump[2]) );
  AOI22_X1 U75 ( .A1(branch_target[2]), .A2(pcsrc), .B1(from_increment_pc[2]), 
        .B2(n15), .ZN(n44) );
endmodule


module writeback ( from_mem_data, from_alu_data, regfile_addr_in, regwrite_in, 
        link, memtoreg, regwrite_out, regfile_data, regfile_addr_out );
  input [31:0] from_mem_data;
  input [31:0] from_alu_data;
  input [4:0] regfile_addr_in;
  output [31:0] regfile_data;
  output [4:0] regfile_addr_out;
  input regwrite_in, link, memtoreg;
  output regwrite_out;
  wire   regwrite_in;
  assign regwrite_out = regwrite_in;

  mux21_NBIT32_1 memtoreg_mux21 ( .A(from_mem_data), .B(from_alu_data), .S(
        memtoreg), .Y(regfile_data) );
  mux21_NBIT5_1 link_mux21 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .B(
        regfile_addr_in), .S(link), .Y(regfile_addr_out) );
endmodule


module MEM_WB_Reg ( clk, rst, controls_in, from_mem_data_in, from_alu_data_in, 
        regfile_addr_in, controls_out, from_mem_data_out, from_alu_data_out, 
        regfile_addr_out );
  input [2:0] controls_in;
  input [31:0] from_mem_data_in;
  input [31:0] from_alu_data_in;
  input [4:0] regfile_addr_in;
  output [2:0] controls_out;
  output [31:0] from_mem_data_out;
  output [31:0] from_alu_data_out;
  output [4:0] regfile_addr_out;
  input clk, rst;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, n74, n81, n82, n83, n84, n85, n86;

  DFF_X1 \regfile_addr_out_reg[4]  ( .D(N74), .CK(clk), .Q(regfile_addr_out[4]) );
  DFF_X1 \regfile_addr_out_reg[3]  ( .D(N73), .CK(clk), .Q(regfile_addr_out[3]) );
  DFF_X1 \regfile_addr_out_reg[2]  ( .D(N72), .CK(clk), .Q(regfile_addr_out[2]) );
  DFF_X1 \regfile_addr_out_reg[1]  ( .D(N71), .CK(clk), .Q(regfile_addr_out[1]) );
  DFF_X1 \regfile_addr_out_reg[0]  ( .D(N70), .CK(clk), .Q(regfile_addr_out[0]) );
  DFF_X1 \controls_out_reg[2]  ( .D(N5), .CK(clk), .Q(controls_out[2]) );
  DFF_X1 \controls_out_reg[1]  ( .D(N4), .CK(clk), .Q(controls_out[1]) );
  DFF_X1 \controls_out_reg[0]  ( .D(N3), .CK(clk), .Q(controls_out[0]) );
  DFF_X1 \from_mem_data_out_reg[31]  ( .D(N37), .CK(clk), .Q(
        from_mem_data_out[31]) );
  DFF_X1 \from_mem_data_out_reg[30]  ( .D(N36), .CK(clk), .Q(
        from_mem_data_out[30]) );
  DFF_X1 \from_mem_data_out_reg[29]  ( .D(N35), .CK(clk), .Q(
        from_mem_data_out[29]) );
  DFF_X1 \from_mem_data_out_reg[28]  ( .D(N34), .CK(clk), .Q(
        from_mem_data_out[28]) );
  DFF_X1 \from_mem_data_out_reg[27]  ( .D(N33), .CK(clk), .Q(
        from_mem_data_out[27]) );
  DFF_X1 \from_mem_data_out_reg[26]  ( .D(N32), .CK(clk), .Q(
        from_mem_data_out[26]) );
  DFF_X1 \from_mem_data_out_reg[25]  ( .D(N31), .CK(clk), .Q(
        from_mem_data_out[25]) );
  DFF_X1 \from_mem_data_out_reg[24]  ( .D(N30), .CK(clk), .Q(
        from_mem_data_out[24]) );
  DFF_X1 \from_mem_data_out_reg[23]  ( .D(N29), .CK(clk), .Q(
        from_mem_data_out[23]) );
  DFF_X1 \from_mem_data_out_reg[22]  ( .D(N28), .CK(clk), .Q(
        from_mem_data_out[22]) );
  DFF_X1 \from_mem_data_out_reg[21]  ( .D(N27), .CK(clk), .Q(
        from_mem_data_out[21]) );
  DFF_X1 \from_mem_data_out_reg[20]  ( .D(N26), .CK(clk), .Q(
        from_mem_data_out[20]) );
  DFF_X1 \from_mem_data_out_reg[19]  ( .D(N25), .CK(clk), .Q(
        from_mem_data_out[19]) );
  DFF_X1 \from_mem_data_out_reg[18]  ( .D(N24), .CK(clk), .Q(
        from_mem_data_out[18]) );
  DFF_X1 \from_mem_data_out_reg[17]  ( .D(N23), .CK(clk), .Q(
        from_mem_data_out[17]) );
  DFF_X1 \from_mem_data_out_reg[16]  ( .D(N22), .CK(clk), .Q(
        from_mem_data_out[16]) );
  DFF_X1 \from_mem_data_out_reg[15]  ( .D(N21), .CK(clk), .Q(
        from_mem_data_out[15]) );
  DFF_X1 \from_mem_data_out_reg[14]  ( .D(N20), .CK(clk), .Q(
        from_mem_data_out[14]) );
  DFF_X1 \from_mem_data_out_reg[13]  ( .D(N19), .CK(clk), .Q(
        from_mem_data_out[13]) );
  DFF_X1 \from_mem_data_out_reg[12]  ( .D(N18), .CK(clk), .Q(
        from_mem_data_out[12]) );
  DFF_X1 \from_mem_data_out_reg[11]  ( .D(N17), .CK(clk), .Q(
        from_mem_data_out[11]) );
  DFF_X1 \from_mem_data_out_reg[10]  ( .D(N16), .CK(clk), .Q(
        from_mem_data_out[10]) );
  DFF_X1 \from_mem_data_out_reg[9]  ( .D(N15), .CK(clk), .Q(
        from_mem_data_out[9]) );
  DFF_X1 \from_mem_data_out_reg[8]  ( .D(N14), .CK(clk), .Q(
        from_mem_data_out[8]) );
  DFF_X1 \from_mem_data_out_reg[7]  ( .D(N13), .CK(clk), .Q(
        from_mem_data_out[7]) );
  DFF_X1 \from_mem_data_out_reg[6]  ( .D(N12), .CK(clk), .Q(
        from_mem_data_out[6]) );
  DFF_X1 \from_mem_data_out_reg[5]  ( .D(N11), .CK(clk), .Q(
        from_mem_data_out[5]) );
  DFF_X1 \from_mem_data_out_reg[4]  ( .D(N10), .CK(clk), .Q(
        from_mem_data_out[4]) );
  DFF_X1 \from_mem_data_out_reg[3]  ( .D(N9), .CK(clk), .Q(
        from_mem_data_out[3]) );
  DFF_X1 \from_mem_data_out_reg[2]  ( .D(N8), .CK(clk), .Q(
        from_mem_data_out[2]) );
  DFF_X1 \from_mem_data_out_reg[1]  ( .D(N7), .CK(clk), .Q(
        from_mem_data_out[1]) );
  DFF_X1 \from_mem_data_out_reg[0]  ( .D(N6), .CK(clk), .Q(
        from_mem_data_out[0]) );
  DFF_X1 \from_alu_data_out_reg[31]  ( .D(N69), .CK(clk), .Q(
        from_alu_data_out[31]) );
  DFF_X1 \from_alu_data_out_reg[30]  ( .D(N68), .CK(clk), .Q(
        from_alu_data_out[30]) );
  DFF_X1 \from_alu_data_out_reg[29]  ( .D(N67), .CK(clk), .Q(
        from_alu_data_out[29]) );
  DFF_X1 \from_alu_data_out_reg[28]  ( .D(N66), .CK(clk), .Q(
        from_alu_data_out[28]) );
  DFF_X1 \from_alu_data_out_reg[27]  ( .D(N65), .CK(clk), .Q(
        from_alu_data_out[27]) );
  DFF_X1 \from_alu_data_out_reg[26]  ( .D(N64), .CK(clk), .Q(
        from_alu_data_out[26]) );
  DFF_X1 \from_alu_data_out_reg[25]  ( .D(N63), .CK(clk), .Q(
        from_alu_data_out[25]) );
  DFF_X1 \from_alu_data_out_reg[24]  ( .D(N62), .CK(clk), .Q(
        from_alu_data_out[24]) );
  DFF_X1 \from_alu_data_out_reg[23]  ( .D(N61), .CK(clk), .Q(
        from_alu_data_out[23]) );
  DFF_X1 \from_alu_data_out_reg[22]  ( .D(N60), .CK(clk), .Q(
        from_alu_data_out[22]) );
  DFF_X1 \from_alu_data_out_reg[21]  ( .D(N59), .CK(clk), .Q(
        from_alu_data_out[21]) );
  DFF_X1 \from_alu_data_out_reg[20]  ( .D(N58), .CK(clk), .Q(
        from_alu_data_out[20]) );
  DFF_X1 \from_alu_data_out_reg[19]  ( .D(N57), .CK(clk), .Q(
        from_alu_data_out[19]) );
  DFF_X1 \from_alu_data_out_reg[18]  ( .D(N56), .CK(clk), .Q(
        from_alu_data_out[18]) );
  DFF_X1 \from_alu_data_out_reg[17]  ( .D(N55), .CK(clk), .Q(
        from_alu_data_out[17]) );
  DFF_X1 \from_alu_data_out_reg[16]  ( .D(N54), .CK(clk), .Q(
        from_alu_data_out[16]) );
  DFF_X1 \from_alu_data_out_reg[15]  ( .D(N53), .CK(clk), .Q(
        from_alu_data_out[15]) );
  DFF_X1 \from_alu_data_out_reg[14]  ( .D(N52), .CK(clk), .Q(
        from_alu_data_out[14]) );
  DFF_X1 \from_alu_data_out_reg[13]  ( .D(N51), .CK(clk), .Q(
        from_alu_data_out[13]) );
  DFF_X1 \from_alu_data_out_reg[12]  ( .D(N50), .CK(clk), .Q(
        from_alu_data_out[12]) );
  DFF_X1 \from_alu_data_out_reg[11]  ( .D(N49), .CK(clk), .Q(
        from_alu_data_out[11]) );
  DFF_X1 \from_alu_data_out_reg[10]  ( .D(N48), .CK(clk), .Q(
        from_alu_data_out[10]) );
  DFF_X1 \from_alu_data_out_reg[9]  ( .D(N47), .CK(clk), .Q(
        from_alu_data_out[9]) );
  DFF_X1 \from_alu_data_out_reg[8]  ( .D(N46), .CK(clk), .Q(
        from_alu_data_out[8]) );
  DFF_X1 \from_alu_data_out_reg[7]  ( .D(N45), .CK(clk), .Q(
        from_alu_data_out[7]) );
  DFF_X1 \from_alu_data_out_reg[6]  ( .D(N44), .CK(clk), .Q(
        from_alu_data_out[6]) );
  DFF_X1 \from_alu_data_out_reg[5]  ( .D(N43), .CK(clk), .Q(
        from_alu_data_out[5]) );
  DFF_X1 \from_alu_data_out_reg[4]  ( .D(N42), .CK(clk), .Q(
        from_alu_data_out[4]) );
  DFF_X1 \from_alu_data_out_reg[3]  ( .D(N41), .CK(clk), .Q(
        from_alu_data_out[3]) );
  DFF_X1 \from_alu_data_out_reg[2]  ( .D(N40), .CK(clk), .Q(
        from_alu_data_out[2]) );
  DFF_X1 \from_alu_data_out_reg[1]  ( .D(N39), .CK(clk), .Q(
        from_alu_data_out[1]) );
  DFF_X1 \from_alu_data_out_reg[0]  ( .D(N38), .CK(clk), .Q(
        from_alu_data_out[0]) );
  BUF_X1 U3 ( .A(n74), .Z(n85) );
  BUF_X1 U4 ( .A(n74), .Z(n81) );
  BUF_X1 U5 ( .A(n74), .Z(n82) );
  BUF_X1 U6 ( .A(n74), .Z(n83) );
  BUF_X1 U7 ( .A(n74), .Z(n84) );
  BUF_X1 U8 ( .A(n74), .Z(n86) );
  AND2_X1 U9 ( .A1(from_mem_data_in[15]), .A2(n81), .ZN(N21) );
  AND2_X1 U10 ( .A1(from_mem_data_in[26]), .A2(n82), .ZN(N32) );
  AND2_X1 U11 ( .A1(from_mem_data_in[23]), .A2(n82), .ZN(N29) );
  AND2_X1 U12 ( .A1(from_mem_data_in[24]), .A2(n82), .ZN(N30) );
  AND2_X1 U13 ( .A1(from_mem_data_in[25]), .A2(n82), .ZN(N31) );
  AND2_X1 U14 ( .A1(from_mem_data_in[27]), .A2(n83), .ZN(N33) );
  AND2_X1 U15 ( .A1(from_mem_data_in[28]), .A2(n83), .ZN(N34) );
  AND2_X1 U16 ( .A1(from_mem_data_in[29]), .A2(n83), .ZN(N35) );
  AND2_X1 U17 ( .A1(from_mem_data_in[30]), .A2(n83), .ZN(N36) );
  AND2_X1 U18 ( .A1(from_mem_data_in[31]), .A2(n83), .ZN(N37) );
  INV_X1 U19 ( .A(rst), .ZN(n74) );
  AND2_X1 U20 ( .A1(from_alu_data_in[0]), .A2(n83), .ZN(N38) );
  AND2_X1 U21 ( .A1(from_alu_data_in[1]), .A2(n83), .ZN(N39) );
  AND2_X1 U22 ( .A1(from_mem_data_in[8]), .A2(n81), .ZN(N14) );
  AND2_X1 U23 ( .A1(from_mem_data_in[9]), .A2(n81), .ZN(N15) );
  AND2_X1 U24 ( .A1(from_mem_data_in[10]), .A2(n81), .ZN(N16) );
  AND2_X1 U25 ( .A1(from_mem_data_in[11]), .A2(n81), .ZN(N17) );
  AND2_X1 U26 ( .A1(from_mem_data_in[12]), .A2(n81), .ZN(N18) );
  AND2_X1 U27 ( .A1(from_mem_data_in[13]), .A2(n81), .ZN(N19) );
  AND2_X1 U28 ( .A1(from_mem_data_in[14]), .A2(n81), .ZN(N20) );
  AND2_X1 U29 ( .A1(from_mem_data_in[7]), .A2(n81), .ZN(N13) );
  AND2_X1 U30 ( .A1(regfile_addr_in[0]), .A2(n86), .ZN(N70) );
  AND2_X1 U31 ( .A1(regfile_addr_in[1]), .A2(n86), .ZN(N71) );
  AND2_X1 U32 ( .A1(regfile_addr_in[2]), .A2(n86), .ZN(N72) );
  AND2_X1 U33 ( .A1(regfile_addr_in[4]), .A2(n86), .ZN(N74) );
  AND2_X1 U34 ( .A1(regfile_addr_in[3]), .A2(n86), .ZN(N73) );
  AND2_X1 U35 ( .A1(from_mem_data_in[16]), .A2(n82), .ZN(N22) );
  AND2_X1 U36 ( .A1(from_mem_data_in[17]), .A2(n82), .ZN(N23) );
  AND2_X1 U37 ( .A1(from_mem_data_in[18]), .A2(n82), .ZN(N24) );
  AND2_X1 U38 ( .A1(from_mem_data_in[19]), .A2(n82), .ZN(N25) );
  AND2_X1 U39 ( .A1(from_mem_data_in[20]), .A2(n82), .ZN(N26) );
  AND2_X1 U40 ( .A1(from_mem_data_in[21]), .A2(n82), .ZN(N27) );
  AND2_X1 U41 ( .A1(from_mem_data_in[22]), .A2(n82), .ZN(N28) );
  AND2_X1 U42 ( .A1(from_alu_data_in[2]), .A2(n83), .ZN(N40) );
  AND2_X1 U43 ( .A1(from_alu_data_in[3]), .A2(n83), .ZN(N41) );
  AND2_X1 U44 ( .A1(from_alu_data_in[4]), .A2(n83), .ZN(N42) );
  AND2_X1 U45 ( .A1(from_alu_data_in[5]), .A2(n83), .ZN(N43) );
  AND2_X1 U46 ( .A1(from_alu_data_in[6]), .A2(n84), .ZN(N44) );
  AND2_X1 U47 ( .A1(from_alu_data_in[7]), .A2(n84), .ZN(N45) );
  AND2_X1 U48 ( .A1(from_alu_data_in[8]), .A2(n84), .ZN(N46) );
  AND2_X1 U49 ( .A1(from_alu_data_in[9]), .A2(n84), .ZN(N47) );
  AND2_X1 U50 ( .A1(from_alu_data_in[10]), .A2(n84), .ZN(N48) );
  AND2_X1 U51 ( .A1(from_alu_data_in[11]), .A2(n84), .ZN(N49) );
  AND2_X1 U52 ( .A1(from_alu_data_in[12]), .A2(n84), .ZN(N50) );
  AND2_X1 U53 ( .A1(from_alu_data_in[13]), .A2(n84), .ZN(N51) );
  AND2_X1 U54 ( .A1(from_alu_data_in[14]), .A2(n84), .ZN(N52) );
  AND2_X1 U55 ( .A1(from_alu_data_in[15]), .A2(n84), .ZN(N53) );
  AND2_X1 U56 ( .A1(from_alu_data_in[16]), .A2(n84), .ZN(N54) );
  AND2_X1 U57 ( .A1(from_alu_data_in[17]), .A2(n85), .ZN(N55) );
  AND2_X1 U58 ( .A1(from_alu_data_in[18]), .A2(n85), .ZN(N56) );
  AND2_X1 U59 ( .A1(from_alu_data_in[19]), .A2(n85), .ZN(N57) );
  AND2_X1 U60 ( .A1(from_alu_data_in[20]), .A2(n85), .ZN(N58) );
  AND2_X1 U61 ( .A1(from_alu_data_in[21]), .A2(n85), .ZN(N59) );
  AND2_X1 U62 ( .A1(from_alu_data_in[22]), .A2(n85), .ZN(N60) );
  AND2_X1 U63 ( .A1(from_alu_data_in[23]), .A2(n85), .ZN(N61) );
  AND2_X1 U64 ( .A1(from_alu_data_in[24]), .A2(n85), .ZN(N62) );
  AND2_X1 U65 ( .A1(from_alu_data_in[25]), .A2(n85), .ZN(N63) );
  AND2_X1 U66 ( .A1(from_alu_data_in[26]), .A2(n85), .ZN(N64) );
  AND2_X1 U67 ( .A1(from_alu_data_in[27]), .A2(n85), .ZN(N65) );
  AND2_X1 U68 ( .A1(from_alu_data_in[28]), .A2(n86), .ZN(N66) );
  AND2_X1 U69 ( .A1(from_alu_data_in[29]), .A2(n86), .ZN(N67) );
  AND2_X1 U70 ( .A1(from_alu_data_in[30]), .A2(n86), .ZN(N68) );
  AND2_X1 U71 ( .A1(from_alu_data_in[31]), .A2(n86), .ZN(N69) );
  AND2_X1 U72 ( .A1(from_mem_data_in[0]), .A2(n85), .ZN(N6) );
  AND2_X1 U73 ( .A1(from_mem_data_in[1]), .A2(n86), .ZN(N7) );
  AND2_X1 U74 ( .A1(from_mem_data_in[2]), .A2(n86), .ZN(N8) );
  AND2_X1 U75 ( .A1(from_mem_data_in[3]), .A2(n86), .ZN(N9) );
  AND2_X1 U76 ( .A1(from_mem_data_in[4]), .A2(n81), .ZN(N10) );
  AND2_X1 U77 ( .A1(from_mem_data_in[5]), .A2(n81), .ZN(N11) );
  AND2_X1 U78 ( .A1(from_mem_data_in[6]), .A2(n81), .ZN(N12) );
  AND2_X1 U79 ( .A1(controls_in[0]), .A2(n82), .ZN(N3) );
  AND2_X1 U80 ( .A1(controls_in[1]), .A2(n83), .ZN(N4) );
  AND2_X1 U81 ( .A1(controls_in[2]), .A2(n84), .ZN(N5) );
endmodule


module memory ( controls_in, PC1_in, PC2_in, takeBranch, addrMem, writeData, 
        RFaddr_in, Data_out_fromRAM, controls_out, dataOut_mem, dataOut_exe, 
        RFaddr_out, unaligned, PCsrc, flush, jump, PC1_out, PC2_out, 
        regwrite_MEM, RFaddr_MEM, forw_addr_MEM, read_op, write_op, nibble, 
        write_byte, Address_toRAM, Data_in );
  input [10:0] controls_in;
  input [31:0] PC1_in;
  input [31:0] PC2_in;
  input [31:0] addrMem;
  input [31:0] writeData;
  input [4:0] RFaddr_in;
  input [31:0] Data_out_fromRAM;
  output [2:0] controls_out;
  output [31:0] dataOut_mem;
  output [31:0] dataOut_exe;
  output [4:0] RFaddr_out;
  output [31:0] PC1_out;
  output [31:0] PC2_out;
  output [4:0] RFaddr_MEM;
  output [31:0] forw_addr_MEM;
  output [1:0] nibble;
  output [31:0] Address_toRAM;
  output [31:0] Data_in;
  input takeBranch;
  output unaligned, PCsrc, flush, jump, regwrite_MEM, read_op, write_op,
         write_byte;
  wire   controls_in_1, controls_in_0, \controls_in[10] , \controls_in[9] ,
         \controls_in[2] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign jump = controls_in_1;
  assign controls_in_1 = controls_in[1];
  assign controls_in_0 = controls_in[0];
  assign controls_out[2] = \controls_in[10] ;
  assign regwrite_MEM = \controls_in[10] ;
  assign \controls_in[10]  = controls_in[10];
  assign controls_out[1] = \controls_in[9] ;
  assign \controls_in[9]  = controls_in[9];
  assign controls_out[0] = \controls_in[2] ;
  assign \controls_in[2]  = controls_in[2];
  assign PC1_out[31] = PC1_in[31];
  assign PC1_out[30] = PC1_in[30];
  assign PC1_out[29] = PC1_in[29];
  assign PC1_out[28] = PC1_in[28];
  assign PC1_out[27] = PC1_in[27];
  assign PC1_out[26] = PC1_in[26];
  assign PC1_out[25] = PC1_in[25];
  assign PC1_out[24] = PC1_in[24];
  assign PC1_out[23] = PC1_in[23];
  assign PC1_out[22] = PC1_in[22];
  assign PC1_out[21] = PC1_in[21];
  assign PC1_out[20] = PC1_in[20];
  assign PC1_out[19] = PC1_in[19];
  assign PC1_out[18] = PC1_in[18];
  assign PC1_out[17] = PC1_in[17];
  assign PC1_out[16] = PC1_in[16];
  assign PC1_out[15] = PC1_in[15];
  assign PC1_out[14] = PC1_in[14];
  assign PC1_out[13] = PC1_in[13];
  assign PC1_out[12] = PC1_in[12];
  assign PC1_out[11] = PC1_in[11];
  assign PC1_out[10] = PC1_in[10];
  assign PC1_out[9] = PC1_in[9];
  assign PC1_out[8] = PC1_in[8];
  assign PC1_out[7] = PC1_in[7];
  assign PC1_out[6] = PC1_in[6];
  assign PC1_out[5] = PC1_in[5];
  assign PC1_out[4] = PC1_in[4];
  assign PC1_out[3] = PC1_in[3];
  assign PC1_out[2] = PC1_in[2];
  assign PC1_out[1] = PC1_in[1];
  assign PC1_out[0] = PC1_in[0];
  assign PC2_out[31] = PC2_in[31];
  assign PC2_out[30] = PC2_in[30];
  assign PC2_out[29] = PC2_in[29];
  assign PC2_out[28] = PC2_in[28];
  assign PC2_out[27] = PC2_in[27];
  assign PC2_out[26] = PC2_in[26];
  assign PC2_out[25] = PC2_in[25];
  assign PC2_out[24] = PC2_in[24];
  assign PC2_out[23] = PC2_in[23];
  assign PC2_out[22] = PC2_in[22];
  assign PC2_out[21] = PC2_in[21];
  assign PC2_out[20] = PC2_in[20];
  assign PC2_out[19] = PC2_in[19];
  assign PC2_out[18] = PC2_in[18];
  assign PC2_out[17] = PC2_in[17];
  assign PC2_out[16] = PC2_in[16];
  assign PC2_out[15] = PC2_in[15];
  assign PC2_out[14] = PC2_in[14];
  assign PC2_out[13] = PC2_in[13];
  assign PC2_out[12] = PC2_in[12];
  assign PC2_out[11] = PC2_in[11];
  assign PC2_out[10] = PC2_in[10];
  assign PC2_out[9] = PC2_in[9];
  assign PC2_out[8] = PC2_in[8];
  assign PC2_out[7] = PC2_in[7];
  assign PC2_out[6] = PC2_in[6];
  assign PC2_out[5] = PC2_in[5];
  assign PC2_out[4] = PC2_in[4];
  assign PC2_out[3] = PC2_in[3];
  assign PC2_out[2] = PC2_in[2];
  assign PC2_out[1] = PC2_in[1];
  assign PC2_out[0] = PC2_in[0];
  assign RFaddr_out[4] = RFaddr_in[4];
  assign RFaddr_MEM[4] = RFaddr_in[4];
  assign RFaddr_out[3] = RFaddr_in[3];
  assign RFaddr_MEM[3] = RFaddr_in[3];
  assign RFaddr_out[2] = RFaddr_in[2];
  assign RFaddr_MEM[2] = RFaddr_in[2];
  assign RFaddr_out[1] = RFaddr_in[1];
  assign RFaddr_MEM[1] = RFaddr_in[1];
  assign RFaddr_out[0] = RFaddr_in[0];
  assign RFaddr_MEM[0] = RFaddr_in[0];
  assign dataOut_exe[31] = addrMem[31];
  assign forw_addr_MEM[31] = addrMem[31];
  assign dataOut_exe[30] = addrMem[30];
  assign forw_addr_MEM[30] = addrMem[30];
  assign dataOut_exe[29] = addrMem[29];
  assign forw_addr_MEM[29] = addrMem[29];
  assign dataOut_exe[28] = addrMem[28];
  assign forw_addr_MEM[28] = addrMem[28];
  assign dataOut_exe[27] = addrMem[27];
  assign forw_addr_MEM[27] = addrMem[27];
  assign dataOut_exe[26] = addrMem[26];
  assign forw_addr_MEM[26] = addrMem[26];
  assign dataOut_exe[25] = addrMem[25];
  assign forw_addr_MEM[25] = addrMem[25];
  assign dataOut_exe[24] = addrMem[24];
  assign forw_addr_MEM[24] = addrMem[24];
  assign dataOut_exe[23] = addrMem[23];
  assign forw_addr_MEM[23] = addrMem[23];
  assign dataOut_exe[22] = addrMem[22];
  assign forw_addr_MEM[22] = addrMem[22];
  assign dataOut_exe[21] = addrMem[21];
  assign forw_addr_MEM[21] = addrMem[21];
  assign dataOut_exe[20] = addrMem[20];
  assign forw_addr_MEM[20] = addrMem[20];
  assign dataOut_exe[19] = addrMem[19];
  assign forw_addr_MEM[19] = addrMem[19];
  assign dataOut_exe[18] = addrMem[18];
  assign forw_addr_MEM[18] = addrMem[18];
  assign dataOut_exe[17] = addrMem[17];
  assign forw_addr_MEM[17] = addrMem[17];
  assign dataOut_exe[16] = addrMem[16];
  assign forw_addr_MEM[16] = addrMem[16];
  assign dataOut_exe[15] = addrMem[15];
  assign forw_addr_MEM[15] = addrMem[15];
  assign dataOut_exe[14] = addrMem[14];
  assign forw_addr_MEM[14] = addrMem[14];
  assign dataOut_exe[13] = addrMem[13];
  assign forw_addr_MEM[13] = addrMem[13];
  assign dataOut_exe[12] = addrMem[12];
  assign forw_addr_MEM[12] = addrMem[12];
  assign dataOut_exe[11] = addrMem[11];
  assign forw_addr_MEM[11] = addrMem[11];
  assign dataOut_exe[10] = addrMem[10];
  assign forw_addr_MEM[10] = addrMem[10];
  assign dataOut_exe[9] = addrMem[9];
  assign forw_addr_MEM[9] = addrMem[9];
  assign dataOut_exe[8] = addrMem[8];
  assign forw_addr_MEM[8] = addrMem[8];
  assign dataOut_exe[7] = addrMem[7];
  assign forw_addr_MEM[7] = addrMem[7];
  assign dataOut_exe[6] = addrMem[6];
  assign forw_addr_MEM[6] = addrMem[6];
  assign dataOut_exe[5] = addrMem[5];
  assign forw_addr_MEM[5] = addrMem[5];
  assign dataOut_exe[4] = addrMem[4];
  assign forw_addr_MEM[4] = addrMem[4];
  assign dataOut_exe[3] = addrMem[3];
  assign forw_addr_MEM[3] = addrMem[3];
  assign dataOut_exe[2] = addrMem[2];
  assign forw_addr_MEM[2] = addrMem[2];
  assign dataOut_exe[1] = addrMem[1];
  assign forw_addr_MEM[1] = addrMem[1];
  assign dataOut_exe[0] = addrMem[0];
  assign forw_addr_MEM[0] = addrMem[0];
  assign Address_toRAM[31] = 1'b0;
  assign Address_toRAM[30] = 1'b0;

  dram_block dram ( .address(addrMem), .data_write(writeData), .mem_op(
        controls_in[8:3]), .Data_out(Data_out_fromRAM), .unaligned(unaligned), 
        .data_read(dataOut_mem), .read_op(read_op), .write_op(write_op), 
        .nibble(nibble), .write_byte(write_byte), .Address_toRAM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, Address_toRAM[29:0]}), .Data_in(Data_in) );
  OR2_X1 U1 ( .A1(PCsrc), .A2(controls_in_1), .ZN(flush) );
  AND2_X1 U2 ( .A1(takeBranch), .A2(controls_in_0), .ZN(PCsrc) );
endmodule


module EX_MEM_Reg ( clk, rst, controls_in, toPC1_in, toPC2_in, takeBranch_in, 
        mem_addr_in, mem_writedata_in, regfile_addr_in, controls_out, 
        toPC1_out, toPC2_out, takeBranch_out, mem_addr_out, mem_writedata_out, 
        regfile_addr_out );
  input [10:0] controls_in;
  input [31:0] toPC1_in;
  input [31:0] toPC2_in;
  input [31:0] mem_addr_in;
  input [31:0] mem_writedata_in;
  input [4:0] regfile_addr_in;
  output [10:0] controls_out;
  output [31:0] toPC1_out;
  output [31:0] toPC2_out;
  output [31:0] mem_addr_out;
  output [31:0] mem_writedata_out;
  output [4:0] regfile_addr_out;
  input clk, rst, takeBranch_in;
  output takeBranch_out;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, n147, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178;

  DFF_X1 \regfile_addr_out_reg[4]  ( .D(N147), .CK(clk), .Q(
        regfile_addr_out[4]) );
  DFF_X1 \regfile_addr_out_reg[3]  ( .D(N146), .CK(clk), .Q(
        regfile_addr_out[3]) );
  DFF_X1 \regfile_addr_out_reg[2]  ( .D(N145), .CK(clk), .Q(
        regfile_addr_out[2]) );
  DFF_X1 \regfile_addr_out_reg[1]  ( .D(N144), .CK(clk), .Q(
        regfile_addr_out[1]) );
  DFF_X1 \regfile_addr_out_reg[0]  ( .D(N143), .CK(clk), .Q(
        regfile_addr_out[0]) );
  DFF_X1 \controls_out_reg[10]  ( .D(N13), .CK(clk), .Q(controls_out[10]) );
  DFF_X1 \controls_out_reg[9]  ( .D(N12), .CK(clk), .Q(controls_out[9]) );
  DFF_X1 \controls_out_reg[8]  ( .D(N11), .CK(clk), .Q(controls_out[8]) );
  DFF_X1 \controls_out_reg[7]  ( .D(N10), .CK(clk), .Q(controls_out[7]) );
  DFF_X1 \controls_out_reg[6]  ( .D(N9), .CK(clk), .Q(controls_out[6]) );
  DFF_X1 \controls_out_reg[5]  ( .D(N8), .CK(clk), .Q(controls_out[5]) );
  DFF_X1 \controls_out_reg[4]  ( .D(N7), .CK(clk), .Q(controls_out[4]) );
  DFF_X1 \controls_out_reg[3]  ( .D(N6), .CK(clk), .Q(controls_out[3]) );
  DFF_X1 \controls_out_reg[2]  ( .D(N5), .CK(clk), .Q(controls_out[2]) );
  DFF_X1 \controls_out_reg[1]  ( .D(N4), .CK(clk), .Q(controls_out[1]) );
  DFF_X1 \controls_out_reg[0]  ( .D(N3), .CK(clk), .Q(controls_out[0]) );
  DFF_X1 \toPC1_out_reg[31]  ( .D(N45), .CK(clk), .Q(toPC1_out[31]) );
  DFF_X1 \toPC1_out_reg[30]  ( .D(N44), .CK(clk), .Q(toPC1_out[30]) );
  DFF_X1 \toPC1_out_reg[29]  ( .D(N43), .CK(clk), .Q(toPC1_out[29]) );
  DFF_X1 \toPC1_out_reg[28]  ( .D(N42), .CK(clk), .Q(toPC1_out[28]) );
  DFF_X1 \toPC1_out_reg[27]  ( .D(N41), .CK(clk), .Q(toPC1_out[27]) );
  DFF_X1 \toPC1_out_reg[26]  ( .D(N40), .CK(clk), .Q(toPC1_out[26]) );
  DFF_X1 \toPC1_out_reg[25]  ( .D(N39), .CK(clk), .Q(toPC1_out[25]) );
  DFF_X1 \toPC1_out_reg[24]  ( .D(N38), .CK(clk), .Q(toPC1_out[24]) );
  DFF_X1 \toPC1_out_reg[23]  ( .D(N37), .CK(clk), .Q(toPC1_out[23]) );
  DFF_X1 \toPC1_out_reg[22]  ( .D(N36), .CK(clk), .Q(toPC1_out[22]) );
  DFF_X1 \toPC1_out_reg[21]  ( .D(N35), .CK(clk), .Q(toPC1_out[21]) );
  DFF_X1 \toPC1_out_reg[20]  ( .D(N34), .CK(clk), .Q(toPC1_out[20]) );
  DFF_X1 \toPC1_out_reg[19]  ( .D(N33), .CK(clk), .Q(toPC1_out[19]) );
  DFF_X1 \toPC1_out_reg[18]  ( .D(N32), .CK(clk), .Q(toPC1_out[18]) );
  DFF_X1 \toPC1_out_reg[17]  ( .D(N31), .CK(clk), .Q(toPC1_out[17]) );
  DFF_X1 \toPC1_out_reg[16]  ( .D(N30), .CK(clk), .Q(toPC1_out[16]) );
  DFF_X1 \toPC1_out_reg[15]  ( .D(N29), .CK(clk), .Q(toPC1_out[15]) );
  DFF_X1 \toPC1_out_reg[14]  ( .D(N28), .CK(clk), .Q(toPC1_out[14]) );
  DFF_X1 \toPC1_out_reg[13]  ( .D(N27), .CK(clk), .Q(toPC1_out[13]) );
  DFF_X1 \toPC1_out_reg[12]  ( .D(N26), .CK(clk), .Q(toPC1_out[12]) );
  DFF_X1 \toPC1_out_reg[11]  ( .D(N25), .CK(clk), .Q(toPC1_out[11]) );
  DFF_X1 \toPC1_out_reg[10]  ( .D(N24), .CK(clk), .Q(toPC1_out[10]) );
  DFF_X1 \toPC1_out_reg[9]  ( .D(N23), .CK(clk), .Q(toPC1_out[9]) );
  DFF_X1 \toPC1_out_reg[8]  ( .D(N22), .CK(clk), .Q(toPC1_out[8]) );
  DFF_X1 \toPC1_out_reg[7]  ( .D(N21), .CK(clk), .Q(toPC1_out[7]) );
  DFF_X1 \toPC1_out_reg[6]  ( .D(N20), .CK(clk), .Q(toPC1_out[6]) );
  DFF_X1 \toPC1_out_reg[5]  ( .D(N19), .CK(clk), .Q(toPC1_out[5]) );
  DFF_X1 \toPC1_out_reg[4]  ( .D(N18), .CK(clk), .Q(toPC1_out[4]) );
  DFF_X1 \toPC1_out_reg[3]  ( .D(N17), .CK(clk), .Q(toPC1_out[3]) );
  DFF_X1 \toPC1_out_reg[2]  ( .D(N16), .CK(clk), .Q(toPC1_out[2]) );
  DFF_X1 \toPC1_out_reg[1]  ( .D(N15), .CK(clk), .Q(toPC1_out[1]) );
  DFF_X1 \toPC1_out_reg[0]  ( .D(N14), .CK(clk), .Q(toPC1_out[0]) );
  DFF_X1 \toPC2_out_reg[31]  ( .D(N77), .CK(clk), .Q(toPC2_out[31]) );
  DFF_X1 \toPC2_out_reg[30]  ( .D(N76), .CK(clk), .Q(toPC2_out[30]) );
  DFF_X1 \toPC2_out_reg[29]  ( .D(N75), .CK(clk), .Q(toPC2_out[29]) );
  DFF_X1 \toPC2_out_reg[28]  ( .D(N74), .CK(clk), .Q(toPC2_out[28]) );
  DFF_X1 \toPC2_out_reg[27]  ( .D(N73), .CK(clk), .Q(toPC2_out[27]) );
  DFF_X1 \toPC2_out_reg[26]  ( .D(N72), .CK(clk), .Q(toPC2_out[26]) );
  DFF_X1 \toPC2_out_reg[25]  ( .D(N71), .CK(clk), .Q(toPC2_out[25]) );
  DFF_X1 \toPC2_out_reg[24]  ( .D(N70), .CK(clk), .Q(toPC2_out[24]) );
  DFF_X1 \toPC2_out_reg[23]  ( .D(N69), .CK(clk), .Q(toPC2_out[23]) );
  DFF_X1 \toPC2_out_reg[22]  ( .D(N68), .CK(clk), .Q(toPC2_out[22]) );
  DFF_X1 \toPC2_out_reg[21]  ( .D(N67), .CK(clk), .Q(toPC2_out[21]) );
  DFF_X1 \toPC2_out_reg[20]  ( .D(N66), .CK(clk), .Q(toPC2_out[20]) );
  DFF_X1 \toPC2_out_reg[19]  ( .D(N65), .CK(clk), .Q(toPC2_out[19]) );
  DFF_X1 \toPC2_out_reg[18]  ( .D(N64), .CK(clk), .Q(toPC2_out[18]) );
  DFF_X1 \toPC2_out_reg[17]  ( .D(N63), .CK(clk), .Q(toPC2_out[17]) );
  DFF_X1 \toPC2_out_reg[16]  ( .D(N62), .CK(clk), .Q(toPC2_out[16]) );
  DFF_X1 \toPC2_out_reg[15]  ( .D(N61), .CK(clk), .Q(toPC2_out[15]) );
  DFF_X1 \toPC2_out_reg[14]  ( .D(N60), .CK(clk), .Q(toPC2_out[14]) );
  DFF_X1 \toPC2_out_reg[13]  ( .D(N59), .CK(clk), .Q(toPC2_out[13]) );
  DFF_X1 \toPC2_out_reg[12]  ( .D(N58), .CK(clk), .Q(toPC2_out[12]) );
  DFF_X1 \toPC2_out_reg[11]  ( .D(N57), .CK(clk), .Q(toPC2_out[11]) );
  DFF_X1 \toPC2_out_reg[10]  ( .D(N56), .CK(clk), .Q(toPC2_out[10]) );
  DFF_X1 \toPC2_out_reg[9]  ( .D(N55), .CK(clk), .Q(toPC2_out[9]) );
  DFF_X1 \toPC2_out_reg[8]  ( .D(N54), .CK(clk), .Q(toPC2_out[8]) );
  DFF_X1 \toPC2_out_reg[7]  ( .D(N53), .CK(clk), .Q(toPC2_out[7]) );
  DFF_X1 \toPC2_out_reg[6]  ( .D(N52), .CK(clk), .Q(toPC2_out[6]) );
  DFF_X1 \toPC2_out_reg[5]  ( .D(N51), .CK(clk), .Q(toPC2_out[5]) );
  DFF_X1 \toPC2_out_reg[4]  ( .D(N50), .CK(clk), .Q(toPC2_out[4]) );
  DFF_X1 \toPC2_out_reg[3]  ( .D(N49), .CK(clk), .Q(toPC2_out[3]) );
  DFF_X1 \toPC2_out_reg[2]  ( .D(N48), .CK(clk), .Q(toPC2_out[2]) );
  DFF_X1 \toPC2_out_reg[1]  ( .D(N47), .CK(clk), .Q(toPC2_out[1]) );
  DFF_X1 \toPC2_out_reg[0]  ( .D(N46), .CK(clk), .Q(toPC2_out[0]) );
  DFF_X1 takeBranch_out_reg ( .D(N78), .CK(clk), .Q(takeBranch_out) );
  DFF_X1 \mem_addr_out_reg[31]  ( .D(N110), .CK(clk), .Q(mem_addr_out[31]) );
  DFF_X1 \mem_addr_out_reg[30]  ( .D(N109), .CK(clk), .Q(mem_addr_out[30]) );
  DFF_X1 \mem_addr_out_reg[29]  ( .D(N108), .CK(clk), .Q(mem_addr_out[29]) );
  DFF_X1 \mem_addr_out_reg[28]  ( .D(N107), .CK(clk), .Q(mem_addr_out[28]) );
  DFF_X1 \mem_addr_out_reg[27]  ( .D(N106), .CK(clk), .Q(mem_addr_out[27]) );
  DFF_X1 \mem_addr_out_reg[26]  ( .D(N105), .CK(clk), .Q(mem_addr_out[26]) );
  DFF_X1 \mem_addr_out_reg[25]  ( .D(N104), .CK(clk), .Q(mem_addr_out[25]) );
  DFF_X1 \mem_addr_out_reg[24]  ( .D(N103), .CK(clk), .Q(mem_addr_out[24]) );
  DFF_X1 \mem_addr_out_reg[23]  ( .D(N102), .CK(clk), .Q(mem_addr_out[23]) );
  DFF_X1 \mem_addr_out_reg[22]  ( .D(N101), .CK(clk), .Q(mem_addr_out[22]) );
  DFF_X1 \mem_addr_out_reg[21]  ( .D(N100), .CK(clk), .Q(mem_addr_out[21]) );
  DFF_X1 \mem_addr_out_reg[20]  ( .D(N99), .CK(clk), .Q(mem_addr_out[20]) );
  DFF_X1 \mem_addr_out_reg[19]  ( .D(N98), .CK(clk), .Q(mem_addr_out[19]) );
  DFF_X1 \mem_addr_out_reg[18]  ( .D(N97), .CK(clk), .Q(mem_addr_out[18]) );
  DFF_X1 \mem_addr_out_reg[17]  ( .D(N96), .CK(clk), .Q(mem_addr_out[17]) );
  DFF_X1 \mem_addr_out_reg[16]  ( .D(N95), .CK(clk), .Q(mem_addr_out[16]) );
  DFF_X1 \mem_addr_out_reg[15]  ( .D(N94), .CK(clk), .Q(mem_addr_out[15]) );
  DFF_X1 \mem_addr_out_reg[14]  ( .D(N93), .CK(clk), .Q(mem_addr_out[14]) );
  DFF_X1 \mem_addr_out_reg[13]  ( .D(N92), .CK(clk), .Q(mem_addr_out[13]) );
  DFF_X1 \mem_addr_out_reg[12]  ( .D(N91), .CK(clk), .Q(mem_addr_out[12]) );
  DFF_X1 \mem_addr_out_reg[11]  ( .D(N90), .CK(clk), .Q(mem_addr_out[11]) );
  DFF_X1 \mem_addr_out_reg[10]  ( .D(N89), .CK(clk), .Q(mem_addr_out[10]) );
  DFF_X1 \mem_addr_out_reg[9]  ( .D(N88), .CK(clk), .Q(mem_addr_out[9]) );
  DFF_X1 \mem_addr_out_reg[8]  ( .D(N87), .CK(clk), .Q(mem_addr_out[8]) );
  DFF_X1 \mem_addr_out_reg[7]  ( .D(N86), .CK(clk), .Q(mem_addr_out[7]) );
  DFF_X1 \mem_addr_out_reg[6]  ( .D(N85), .CK(clk), .Q(mem_addr_out[6]) );
  DFF_X1 \mem_addr_out_reg[5]  ( .D(N84), .CK(clk), .Q(mem_addr_out[5]) );
  DFF_X1 \mem_addr_out_reg[4]  ( .D(N83), .CK(clk), .Q(mem_addr_out[4]) );
  DFF_X1 \mem_addr_out_reg[3]  ( .D(N82), .CK(clk), .Q(mem_addr_out[3]) );
  DFF_X1 \mem_addr_out_reg[2]  ( .D(N81), .CK(clk), .Q(mem_addr_out[2]) );
  DFF_X1 \mem_addr_out_reg[1]  ( .D(N80), .CK(clk), .Q(mem_addr_out[1]) );
  DFF_X1 \mem_addr_out_reg[0]  ( .D(N79), .CK(clk), .Q(mem_addr_out[0]) );
  DFF_X1 \mem_writedata_out_reg[31]  ( .D(N142), .CK(clk), .Q(
        mem_writedata_out[31]) );
  DFF_X1 \mem_writedata_out_reg[30]  ( .D(N141), .CK(clk), .Q(
        mem_writedata_out[30]) );
  DFF_X1 \mem_writedata_out_reg[29]  ( .D(N140), .CK(clk), .Q(
        mem_writedata_out[29]) );
  DFF_X1 \mem_writedata_out_reg[28]  ( .D(N139), .CK(clk), .Q(
        mem_writedata_out[28]) );
  DFF_X1 \mem_writedata_out_reg[27]  ( .D(N138), .CK(clk), .Q(
        mem_writedata_out[27]) );
  DFF_X1 \mem_writedata_out_reg[26]  ( .D(N137), .CK(clk), .Q(
        mem_writedata_out[26]) );
  DFF_X1 \mem_writedata_out_reg[25]  ( .D(N136), .CK(clk), .Q(
        mem_writedata_out[25]) );
  DFF_X1 \mem_writedata_out_reg[24]  ( .D(N135), .CK(clk), .Q(
        mem_writedata_out[24]) );
  DFF_X1 \mem_writedata_out_reg[23]  ( .D(N134), .CK(clk), .Q(
        mem_writedata_out[23]) );
  DFF_X1 \mem_writedata_out_reg[22]  ( .D(N133), .CK(clk), .Q(
        mem_writedata_out[22]) );
  DFF_X1 \mem_writedata_out_reg[21]  ( .D(N132), .CK(clk), .Q(
        mem_writedata_out[21]) );
  DFF_X1 \mem_writedata_out_reg[20]  ( .D(N131), .CK(clk), .Q(
        mem_writedata_out[20]) );
  DFF_X1 \mem_writedata_out_reg[19]  ( .D(N130), .CK(clk), .Q(
        mem_writedata_out[19]) );
  DFF_X1 \mem_writedata_out_reg[18]  ( .D(N129), .CK(clk), .Q(
        mem_writedata_out[18]) );
  DFF_X1 \mem_writedata_out_reg[17]  ( .D(N128), .CK(clk), .Q(
        mem_writedata_out[17]) );
  DFF_X1 \mem_writedata_out_reg[16]  ( .D(N127), .CK(clk), .Q(
        mem_writedata_out[16]) );
  DFF_X1 \mem_writedata_out_reg[15]  ( .D(N126), .CK(clk), .Q(
        mem_writedata_out[15]) );
  DFF_X1 \mem_writedata_out_reg[14]  ( .D(N125), .CK(clk), .Q(
        mem_writedata_out[14]) );
  DFF_X1 \mem_writedata_out_reg[13]  ( .D(N124), .CK(clk), .Q(
        mem_writedata_out[13]) );
  DFF_X1 \mem_writedata_out_reg[12]  ( .D(N123), .CK(clk), .Q(
        mem_writedata_out[12]) );
  DFF_X1 \mem_writedata_out_reg[11]  ( .D(N122), .CK(clk), .Q(
        mem_writedata_out[11]) );
  DFF_X1 \mem_writedata_out_reg[10]  ( .D(N121), .CK(clk), .Q(
        mem_writedata_out[10]) );
  DFF_X1 \mem_writedata_out_reg[9]  ( .D(N120), .CK(clk), .Q(
        mem_writedata_out[9]) );
  DFF_X1 \mem_writedata_out_reg[8]  ( .D(N119), .CK(clk), .Q(
        mem_writedata_out[8]) );
  DFF_X1 \mem_writedata_out_reg[7]  ( .D(N118), .CK(clk), .Q(
        mem_writedata_out[7]) );
  DFF_X1 \mem_writedata_out_reg[6]  ( .D(N117), .CK(clk), .Q(
        mem_writedata_out[6]) );
  DFF_X1 \mem_writedata_out_reg[5]  ( .D(N116), .CK(clk), .Q(
        mem_writedata_out[5]) );
  DFF_X1 \mem_writedata_out_reg[4]  ( .D(N115), .CK(clk), .Q(
        mem_writedata_out[4]) );
  DFF_X1 \mem_writedata_out_reg[3]  ( .D(N114), .CK(clk), .Q(
        mem_writedata_out[3]) );
  DFF_X1 \mem_writedata_out_reg[2]  ( .D(N113), .CK(clk), .Q(
        mem_writedata_out[2]) );
  DFF_X1 \mem_writedata_out_reg[1]  ( .D(N112), .CK(clk), .Q(
        mem_writedata_out[1]) );
  DFF_X1 \mem_writedata_out_reg[0]  ( .D(N111), .CK(clk), .Q(
        mem_writedata_out[0]) );
  BUF_X1 U3 ( .A(n166), .Z(n177) );
  BUF_X1 U4 ( .A(n164), .Z(n170) );
  BUF_X1 U5 ( .A(n165), .Z(n172) );
  BUF_X1 U6 ( .A(n165), .Z(n173) );
  BUF_X1 U7 ( .A(n165), .Z(n174) );
  BUF_X1 U8 ( .A(n165), .Z(n175) );
  BUF_X1 U9 ( .A(n165), .Z(n176) );
  BUF_X1 U10 ( .A(n164), .Z(n167) );
  BUF_X1 U11 ( .A(n164), .Z(n168) );
  BUF_X1 U12 ( .A(n164), .Z(n169) );
  BUF_X1 U13 ( .A(n164), .Z(n171) );
  BUF_X1 U14 ( .A(n166), .Z(n178) );
  BUF_X1 U15 ( .A(n147), .Z(n165) );
  BUF_X1 U16 ( .A(n147), .Z(n164) );
  BUF_X1 U17 ( .A(n147), .Z(n166) );
  AND2_X1 U18 ( .A1(takeBranch_in), .A2(n177), .ZN(N78) );
  INV_X1 U19 ( .A(rst), .ZN(n147) );
  AND2_X1 U20 ( .A1(mem_writedata_in[0]), .A2(n168), .ZN(N111) );
  AND2_X1 U21 ( .A1(mem_writedata_in[1]), .A2(n168), .ZN(N112) );
  AND2_X1 U22 ( .A1(mem_writedata_in[2]), .A2(n168), .ZN(N113) );
  AND2_X1 U23 ( .A1(mem_writedata_in[3]), .A2(n168), .ZN(N114) );
  AND2_X1 U24 ( .A1(mem_writedata_in[4]), .A2(n168), .ZN(N115) );
  AND2_X1 U25 ( .A1(mem_writedata_in[5]), .A2(n168), .ZN(N116) );
  AND2_X1 U26 ( .A1(mem_writedata_in[6]), .A2(n168), .ZN(N117) );
  AND2_X1 U27 ( .A1(mem_writedata_in[7]), .A2(n168), .ZN(N118) );
  AND2_X1 U28 ( .A1(mem_writedata_in[8]), .A2(n168), .ZN(N119) );
  AND2_X1 U29 ( .A1(mem_writedata_in[9]), .A2(n168), .ZN(N120) );
  AND2_X1 U30 ( .A1(mem_writedata_in[10]), .A2(n169), .ZN(N121) );
  AND2_X1 U31 ( .A1(mem_writedata_in[11]), .A2(n169), .ZN(N122) );
  AND2_X1 U32 ( .A1(mem_writedata_in[12]), .A2(n169), .ZN(N123) );
  AND2_X1 U33 ( .A1(mem_writedata_in[13]), .A2(n169), .ZN(N124) );
  AND2_X1 U34 ( .A1(mem_writedata_in[14]), .A2(n169), .ZN(N125) );
  AND2_X1 U35 ( .A1(mem_writedata_in[15]), .A2(n169), .ZN(N126) );
  AND2_X1 U36 ( .A1(mem_writedata_in[16]), .A2(n169), .ZN(N127) );
  AND2_X1 U37 ( .A1(mem_writedata_in[17]), .A2(n169), .ZN(N128) );
  AND2_X1 U38 ( .A1(mem_writedata_in[18]), .A2(n169), .ZN(N129) );
  AND2_X1 U39 ( .A1(mem_writedata_in[19]), .A2(n169), .ZN(N130) );
  AND2_X1 U40 ( .A1(mem_writedata_in[20]), .A2(n169), .ZN(N131) );
  AND2_X1 U41 ( .A1(mem_writedata_in[21]), .A2(n170), .ZN(N132) );
  AND2_X1 U42 ( .A1(mem_writedata_in[22]), .A2(n170), .ZN(N133) );
  AND2_X1 U43 ( .A1(mem_writedata_in[23]), .A2(n170), .ZN(N134) );
  AND2_X1 U44 ( .A1(mem_writedata_in[24]), .A2(n170), .ZN(N135) );
  AND2_X1 U45 ( .A1(mem_writedata_in[25]), .A2(n170), .ZN(N136) );
  AND2_X1 U46 ( .A1(mem_writedata_in[26]), .A2(n170), .ZN(N137) );
  AND2_X1 U47 ( .A1(mem_writedata_in[27]), .A2(n170), .ZN(N138) );
  AND2_X1 U48 ( .A1(mem_writedata_in[28]), .A2(n170), .ZN(N139) );
  AND2_X1 U49 ( .A1(mem_writedata_in[29]), .A2(n170), .ZN(N140) );
  AND2_X1 U50 ( .A1(mem_writedata_in[30]), .A2(n170), .ZN(N141) );
  AND2_X1 U51 ( .A1(mem_writedata_in[31]), .A2(n170), .ZN(N142) );
  AND2_X1 U52 ( .A1(mem_addr_in[0]), .A2(n177), .ZN(N79) );
  AND2_X1 U53 ( .A1(mem_addr_in[1]), .A2(n177), .ZN(N80) );
  AND2_X1 U54 ( .A1(mem_addr_in[2]), .A2(n177), .ZN(N81) );
  AND2_X1 U55 ( .A1(mem_addr_in[3]), .A2(n177), .ZN(N82) );
  AND2_X1 U56 ( .A1(mem_addr_in[4]), .A2(n177), .ZN(N83) );
  AND2_X1 U57 ( .A1(mem_addr_in[5]), .A2(n177), .ZN(N84) );
  AND2_X1 U58 ( .A1(mem_addr_in[6]), .A2(n177), .ZN(N85) );
  AND2_X1 U59 ( .A1(mem_addr_in[7]), .A2(n177), .ZN(N86) );
  AND2_X1 U60 ( .A1(mem_addr_in[8]), .A2(n177), .ZN(N87) );
  AND2_X1 U61 ( .A1(mem_addr_in[21]), .A2(n167), .ZN(N100) );
  AND2_X1 U62 ( .A1(mem_addr_in[22]), .A2(n167), .ZN(N101) );
  AND2_X1 U63 ( .A1(mem_addr_in[23]), .A2(n167), .ZN(N102) );
  AND2_X1 U64 ( .A1(mem_addr_in[24]), .A2(n167), .ZN(N103) );
  AND2_X1 U65 ( .A1(mem_addr_in[25]), .A2(n167), .ZN(N104) );
  AND2_X1 U66 ( .A1(mem_addr_in[26]), .A2(n167), .ZN(N105) );
  AND2_X1 U67 ( .A1(mem_addr_in[27]), .A2(n167), .ZN(N106) );
  AND2_X1 U68 ( .A1(mem_addr_in[28]), .A2(n167), .ZN(N107) );
  AND2_X1 U69 ( .A1(mem_addr_in[29]), .A2(n167), .ZN(N108) );
  AND2_X1 U70 ( .A1(mem_addr_in[30]), .A2(n167), .ZN(N109) );
  AND2_X1 U71 ( .A1(mem_addr_in[31]), .A2(n168), .ZN(N110) );
  AND2_X1 U72 ( .A1(toPC2_in[0]), .A2(n174), .ZN(N46) );
  AND2_X1 U73 ( .A1(toPC2_in[1]), .A2(n174), .ZN(N47) );
  AND2_X1 U74 ( .A1(toPC2_in[2]), .A2(n174), .ZN(N48) );
  AND2_X1 U75 ( .A1(toPC2_in[3]), .A2(n174), .ZN(N49) );
  AND2_X1 U76 ( .A1(toPC2_in[4]), .A2(n174), .ZN(N50) );
  AND2_X1 U77 ( .A1(toPC2_in[5]), .A2(n174), .ZN(N51) );
  AND2_X1 U78 ( .A1(toPC2_in[6]), .A2(n174), .ZN(N52) );
  AND2_X1 U79 ( .A1(toPC2_in[7]), .A2(n174), .ZN(N53) );
  AND2_X1 U80 ( .A1(toPC2_in[8]), .A2(n174), .ZN(N54) );
  AND2_X1 U81 ( .A1(toPC2_in[9]), .A2(n175), .ZN(N55) );
  AND2_X1 U82 ( .A1(toPC2_in[10]), .A2(n175), .ZN(N56) );
  AND2_X1 U83 ( .A1(toPC2_in[11]), .A2(n175), .ZN(N57) );
  AND2_X1 U84 ( .A1(toPC2_in[12]), .A2(n175), .ZN(N58) );
  AND2_X1 U85 ( .A1(toPC2_in[13]), .A2(n175), .ZN(N59) );
  AND2_X1 U86 ( .A1(toPC2_in[14]), .A2(n175), .ZN(N60) );
  AND2_X1 U87 ( .A1(toPC2_in[15]), .A2(n175), .ZN(N61) );
  AND2_X1 U88 ( .A1(toPC2_in[16]), .A2(n175), .ZN(N62) );
  AND2_X1 U89 ( .A1(toPC2_in[17]), .A2(n175), .ZN(N63) );
  AND2_X1 U90 ( .A1(toPC2_in[18]), .A2(n175), .ZN(N64) );
  AND2_X1 U91 ( .A1(toPC2_in[19]), .A2(n175), .ZN(N65) );
  AND2_X1 U92 ( .A1(toPC2_in[20]), .A2(n176), .ZN(N66) );
  AND2_X1 U93 ( .A1(toPC2_in[21]), .A2(n176), .ZN(N67) );
  AND2_X1 U94 ( .A1(toPC2_in[22]), .A2(n176), .ZN(N68) );
  AND2_X1 U95 ( .A1(toPC2_in[23]), .A2(n176), .ZN(N69) );
  AND2_X1 U96 ( .A1(toPC2_in[24]), .A2(n176), .ZN(N70) );
  AND2_X1 U97 ( .A1(toPC2_in[25]), .A2(n176), .ZN(N71) );
  AND2_X1 U98 ( .A1(toPC2_in[26]), .A2(n176), .ZN(N72) );
  AND2_X1 U99 ( .A1(toPC2_in[27]), .A2(n176), .ZN(N73) );
  AND2_X1 U100 ( .A1(toPC2_in[28]), .A2(n176), .ZN(N74) );
  AND2_X1 U101 ( .A1(toPC2_in[29]), .A2(n176), .ZN(N75) );
  AND2_X1 U102 ( .A1(toPC2_in[30]), .A2(n176), .ZN(N76) );
  AND2_X1 U103 ( .A1(toPC2_in[31]), .A2(n177), .ZN(N77) );
  AND2_X1 U104 ( .A1(toPC1_in[0]), .A2(n170), .ZN(N14) );
  AND2_X1 U105 ( .A1(toPC1_in[1]), .A2(n171), .ZN(N15) );
  AND2_X1 U106 ( .A1(toPC1_in[2]), .A2(n171), .ZN(N16) );
  AND2_X1 U107 ( .A1(toPC1_in[3]), .A2(n171), .ZN(N17) );
  AND2_X1 U108 ( .A1(toPC1_in[4]), .A2(n171), .ZN(N18) );
  AND2_X1 U109 ( .A1(toPC1_in[5]), .A2(n171), .ZN(N19) );
  AND2_X1 U110 ( .A1(toPC1_in[6]), .A2(n171), .ZN(N20) );
  AND2_X1 U111 ( .A1(toPC1_in[7]), .A2(n171), .ZN(N21) );
  AND2_X1 U112 ( .A1(toPC1_in[8]), .A2(n172), .ZN(N22) );
  AND2_X1 U113 ( .A1(toPC1_in[9]), .A2(n172), .ZN(N23) );
  AND2_X1 U114 ( .A1(toPC1_in[10]), .A2(n172), .ZN(N24) );
  AND2_X1 U115 ( .A1(toPC1_in[11]), .A2(n172), .ZN(N25) );
  AND2_X1 U116 ( .A1(toPC1_in[12]), .A2(n172), .ZN(N26) );
  AND2_X1 U117 ( .A1(toPC1_in[13]), .A2(n172), .ZN(N27) );
  AND2_X1 U118 ( .A1(toPC1_in[14]), .A2(n172), .ZN(N28) );
  AND2_X1 U119 ( .A1(toPC1_in[15]), .A2(n172), .ZN(N29) );
  AND2_X1 U120 ( .A1(toPC1_in[16]), .A2(n172), .ZN(N30) );
  AND2_X1 U121 ( .A1(toPC1_in[17]), .A2(n172), .ZN(N31) );
  AND2_X1 U122 ( .A1(toPC1_in[18]), .A2(n172), .ZN(N32) );
  AND2_X1 U123 ( .A1(toPC1_in[19]), .A2(n173), .ZN(N33) );
  AND2_X1 U124 ( .A1(toPC1_in[20]), .A2(n173), .ZN(N34) );
  AND2_X1 U125 ( .A1(toPC1_in[21]), .A2(n173), .ZN(N35) );
  AND2_X1 U126 ( .A1(toPC1_in[22]), .A2(n173), .ZN(N36) );
  AND2_X1 U127 ( .A1(toPC1_in[23]), .A2(n173), .ZN(N37) );
  AND2_X1 U128 ( .A1(toPC1_in[24]), .A2(n173), .ZN(N38) );
  AND2_X1 U129 ( .A1(toPC1_in[25]), .A2(n173), .ZN(N39) );
  AND2_X1 U130 ( .A1(toPC1_in[26]), .A2(n173), .ZN(N40) );
  AND2_X1 U131 ( .A1(toPC1_in[27]), .A2(n173), .ZN(N41) );
  AND2_X1 U132 ( .A1(toPC1_in[28]), .A2(n173), .ZN(N42) );
  AND2_X1 U133 ( .A1(toPC1_in[29]), .A2(n173), .ZN(N43) );
  AND2_X1 U134 ( .A1(toPC1_in[30]), .A2(n174), .ZN(N44) );
  AND2_X1 U135 ( .A1(toPC1_in[31]), .A2(n174), .ZN(N45) );
  AND2_X1 U136 ( .A1(controls_in[0]), .A2(n172), .ZN(N3) );
  AND2_X1 U137 ( .A1(controls_in[1]), .A2(n173), .ZN(N4) );
  AND2_X1 U138 ( .A1(controls_in[2]), .A2(n174), .ZN(N5) );
  AND2_X1 U139 ( .A1(controls_in[3]), .A2(n175), .ZN(N6) );
  AND2_X1 U140 ( .A1(controls_in[4]), .A2(n176), .ZN(N7) );
  AND2_X1 U141 ( .A1(controls_in[5]), .A2(n177), .ZN(N8) );
  AND2_X1 U142 ( .A1(controls_in[7]), .A2(n167), .ZN(N10) );
  AND2_X1 U143 ( .A1(controls_in[8]), .A2(n167), .ZN(N11) );
  AND2_X1 U144 ( .A1(controls_in[9]), .A2(n168), .ZN(N12) );
  AND2_X1 U145 ( .A1(controls_in[10]), .A2(n169), .ZN(N13) );
  AND2_X1 U146 ( .A1(regfile_addr_in[0]), .A2(n171), .ZN(N143) );
  AND2_X1 U147 ( .A1(regfile_addr_in[1]), .A2(n171), .ZN(N144) );
  AND2_X1 U148 ( .A1(regfile_addr_in[2]), .A2(n171), .ZN(N145) );
  AND2_X1 U149 ( .A1(regfile_addr_in[3]), .A2(n171), .ZN(N146) );
  AND2_X1 U150 ( .A1(regfile_addr_in[4]), .A2(n171), .ZN(N147) );
  AND2_X1 U151 ( .A1(mem_addr_in[9]), .A2(n178), .ZN(N88) );
  AND2_X1 U152 ( .A1(mem_addr_in[10]), .A2(n178), .ZN(N89) );
  AND2_X1 U153 ( .A1(mem_addr_in[11]), .A2(n178), .ZN(N90) );
  AND2_X1 U154 ( .A1(mem_addr_in[12]), .A2(n178), .ZN(N91) );
  AND2_X1 U155 ( .A1(mem_addr_in[13]), .A2(n178), .ZN(N92) );
  AND2_X1 U156 ( .A1(mem_addr_in[14]), .A2(n178), .ZN(N93) );
  AND2_X1 U157 ( .A1(mem_addr_in[15]), .A2(n178), .ZN(N94) );
  AND2_X1 U158 ( .A1(mem_addr_in[16]), .A2(n178), .ZN(N95) );
  AND2_X1 U159 ( .A1(mem_addr_in[17]), .A2(n178), .ZN(N96) );
  AND2_X1 U160 ( .A1(mem_addr_in[18]), .A2(n178), .ZN(N97) );
  AND2_X1 U161 ( .A1(mem_addr_in[19]), .A2(n178), .ZN(N98) );
  AND2_X1 U162 ( .A1(controls_in[6]), .A2(n178), .ZN(N9) );
  AND2_X1 U163 ( .A1(mem_addr_in[20]), .A2(n166), .ZN(N99) );
endmodule


module execute ( clk, rst, controls_in, ext25_0, nextPC, op_A, op_B, ext15_0, 
        inst15_0, rt_inst, rd_inst, rs_inst, unaligned, forw_dataWB, 
        forw_dataMEM, RFaddr_WB, RFaddr_MEM, regwriteWB, regwriteMEM, 
        controls_out, toPC1, toPC2, branchTaken, addrMem, writeData, addrRF, 
        IDEX_rt, IDEX_memread );
  input [21:0] controls_in;
  input [31:0] ext25_0;
  input [31:0] nextPC;
  input [31:0] op_A;
  input [31:0] op_B;
  input [31:0] ext15_0;
  input [15:0] inst15_0;
  input [4:0] rt_inst;
  input [4:0] rd_inst;
  input [4:0] rs_inst;
  input [31:0] forw_dataWB;
  input [31:0] forw_dataMEM;
  input [4:0] RFaddr_WB;
  input [4:0] RFaddr_MEM;
  output [10:0] controls_out;
  output [31:0] toPC1;
  output [31:0] toPC2;
  output [31:0] addrMem;
  output [31:0] writeData;
  output [4:0] addrRF;
  output [4:0] IDEX_rt;
  output [3:0] IDEX_memread;
  input clk, rst, unaligned, regwriteWB, regwriteMEM;
  output branchTaken;
  wire   controls_in_20, controls_in_19, controls_in_17, controls_in_16,
         controls_in_15, controls_in_14, \controls_in[21] , \controls_in[18] ,
         \controls_in[13] , \controls_in[12] , \controls_in[11] ,
         \controls_in[10] , \controls_in[9] , \controls_in[8] ,
         \controls_in[7] , \controls_in[6] , \controls_in[5] , zero_i, ovf_i,
         \resAdd1_i[9] , \resAdd1_i[8] , \resAdd1_i[7] , \resAdd1_i[6] ,
         \resAdd1_i[5] , \resAdd1_i[4] , \resAdd1_i[3] , \resAdd1_i[31] ,
         \resAdd1_i[30] , \resAdd1_i[2] , \resAdd1_i[29] , \resAdd1_i[28] ,
         \resAdd1_i[27] , \resAdd1_i[26] , \resAdd1_i[25] , \resAdd1_i[24] ,
         \resAdd1_i[23] , \resAdd1_i[22] , \resAdd1_i[21] , \resAdd1_i[20] ,
         \resAdd1_i[1] , \resAdd1_i[19] , \resAdd1_i[18] , \resAdd1_i[17] ,
         \resAdd1_i[16] , \resAdd1_i[15] , \resAdd1_i[14] , \resAdd1_i[13] ,
         \resAdd1_i[12] , \resAdd1_i[11] , \resAdd1_i[10] , \resAdd1_i[0] ,
         \link_value_i[9] , \link_value_i[8] , \link_value_i[7] ,
         \link_value_i[6] , \link_value_i[5] , \link_value_i[4] ,
         \link_value_i[3] , \link_value_i[31] , \link_value_i[30] ,
         \link_value_i[2] , \link_value_i[29] , \link_value_i[28] ,
         \link_value_i[27] , \link_value_i[26] , \link_value_i[25] ,
         \link_value_i[24] , \link_value_i[23] , \link_value_i[22] ,
         \link_value_i[21] , \link_value_i[20] , \link_value_i[1] ,
         \link_value_i[19] , \link_value_i[18] , \link_value_i[17] ,
         \link_value_i[16] , \link_value_i[15] , \link_value_i[14] ,
         \link_value_i[13] , \link_value_i[12] , \link_value_i[11] ,
         \link_value_i[10] , \link_value_i[0] , \link2lhi_wire_i[9] ,
         \link2lhi_wire_i[8] , \link2lhi_wire_i[7] , \link2lhi_wire_i[6] ,
         \link2lhi_wire_i[5] , \link2lhi_wire_i[4] , \link2lhi_wire_i[3] ,
         \link2lhi_wire_i[31] , \link2lhi_wire_i[30] , \link2lhi_wire_i[2] ,
         \link2lhi_wire_i[29] , \link2lhi_wire_i[28] , \link2lhi_wire_i[27] ,
         \link2lhi_wire_i[26] , \link2lhi_wire_i[25] , \link2lhi_wire_i[24] ,
         \link2lhi_wire_i[23] , \link2lhi_wire_i[22] , \link2lhi_wire_i[21] ,
         \link2lhi_wire_i[20] , \link2lhi_wire_i[1] , \link2lhi_wire_i[19] ,
         \link2lhi_wire_i[18] , \link2lhi_wire_i[17] , \link2lhi_wire_i[16] ,
         \link2lhi_wire_i[15] , \link2lhi_wire_i[14] , \link2lhi_wire_i[13] ,
         \link2lhi_wire_i[12] , \link2lhi_wire_i[11] , \link2lhi_wire_i[10] ,
         \link2lhi_wire_i[0] , \lhi2mov_wire_i[9] , \lhi2mov_wire_i[8] ,
         \lhi2mov_wire_i[7] , \lhi2mov_wire_i[6] , \lhi2mov_wire_i[5] ,
         \lhi2mov_wire_i[4] , \lhi2mov_wire_i[3] , \lhi2mov_wire_i[31] ,
         \lhi2mov_wire_i[30] , \lhi2mov_wire_i[2] , \lhi2mov_wire_i[29] ,
         \lhi2mov_wire_i[28] , \lhi2mov_wire_i[27] , \lhi2mov_wire_i[26] ,
         \lhi2mov_wire_i[25] , \lhi2mov_wire_i[24] , \lhi2mov_wire_i[23] ,
         \lhi2mov_wire_i[22] , \lhi2mov_wire_i[21] , \lhi2mov_wire_i[20] ,
         \lhi2mov_wire_i[1] , \lhi2mov_wire_i[19] , \lhi2mov_wire_i[18] ,
         \lhi2mov_wire_i[17] , \lhi2mov_wire_i[16] , \lhi2mov_wire_i[15] ,
         \lhi2mov_wire_i[14] , \lhi2mov_wire_i[13] , \lhi2mov_wire_i[12] ,
         \lhi2mov_wire_i[11] , \lhi2mov_wire_i[10] , \lhi2mov_wire_i[0] ;
  wire   [31:0] A_inALU_i;
  wire   [31:0] res_outALU_i;
  wire   [31:0] lhi_value_i;
  wire   [31:0] psw_status_i;
  wire   [31:0] B_inALU_i;
  wire   [1:0] forwardA_i;
  wire   [1:0] forwardB_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45;
  assign controls_in_20 = controls_in[20];
  assign controls_in_19 = controls_in[19];
  assign controls_in_17 = controls_in[17];
  assign controls_in_16 = controls_in[16];
  assign controls_in_15 = controls_in[15];
  assign controls_in_14 = controls_in[14];
  assign controls_out[10] = \controls_in[21] ;
  assign \controls_in[21]  = controls_in[21];
  assign controls_out[9] = \controls_in[18] ;
  assign \controls_in[18]  = controls_in[18];
  assign controls_out[8] = \controls_in[13] ;
  assign \controls_in[13]  = controls_in[13];
  assign controls_out[7] = \controls_in[12] ;
  assign \controls_in[12]  = controls_in[12];
  assign controls_out[6] = \controls_in[11] ;
  assign IDEX_memread[3] = \controls_in[11] ;
  assign \controls_in[11]  = controls_in[11];
  assign controls_out[5] = \controls_in[10] ;
  assign IDEX_memread[2] = \controls_in[10] ;
  assign \controls_in[10]  = controls_in[10];
  assign controls_out[4] = \controls_in[9] ;
  assign IDEX_memread[1] = \controls_in[9] ;
  assign \controls_in[9]  = controls_in[9];
  assign controls_out[3] = \controls_in[8] ;
  assign IDEX_memread[0] = \controls_in[8] ;
  assign \controls_in[8]  = controls_in[8];
  assign controls_out[2] = \controls_in[7] ;
  assign \controls_in[7]  = controls_in[7];
  assign controls_out[1] = \controls_in[6] ;
  assign \controls_in[6]  = controls_in[6];
  assign controls_out[0] = \controls_in[5] ;
  assign \controls_in[5]  = controls_in[5];
  assign IDEX_rt[4] = rt_inst[4];
  assign IDEX_rt[3] = rt_inst[3];
  assign IDEX_rt[2] = rt_inst[2];
  assign IDEX_rt[1] = rt_inst[1];
  assign IDEX_rt[0] = rt_inst[0];

  adder_0 adder1 ( .a(ext25_0), .b(nextPC), .res({\resAdd1_i[31] , 
        \resAdd1_i[30] , \resAdd1_i[29] , \resAdd1_i[28] , \resAdd1_i[27] , 
        \resAdd1_i[26] , \resAdd1_i[25] , \resAdd1_i[24] , \resAdd1_i[23] , 
        \resAdd1_i[22] , \resAdd1_i[21] , \resAdd1_i[20] , \resAdd1_i[19] , 
        \resAdd1_i[18] , \resAdd1_i[17] , \resAdd1_i[16] , \resAdd1_i[15] , 
        \resAdd1_i[14] , \resAdd1_i[13] , \resAdd1_i[12] , \resAdd1_i[11] , 
        \resAdd1_i[10] , \resAdd1_i[9] , \resAdd1_i[8] , \resAdd1_i[7] , 
        \resAdd1_i[6] , \resAdd1_i[5] , \resAdd1_i[4] , \resAdd1_i[3] , 
        \resAdd1_i[2] , \resAdd1_i[1] , \resAdd1_i[0] }) );
  adder_2 adder2 ( .a(nextPC), .b(ext15_0), .res(toPC2) );
  adder_1 plus4_adder ( .a(nextPC), .b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .res({\link_value_i[31] , \link_value_i[30] , 
        \link_value_i[29] , \link_value_i[28] , \link_value_i[27] , 
        \link_value_i[26] , \link_value_i[25] , \link_value_i[24] , 
        \link_value_i[23] , \link_value_i[22] , \link_value_i[21] , 
        \link_value_i[20] , \link_value_i[19] , \link_value_i[18] , 
        \link_value_i[17] , \link_value_i[16] , \link_value_i[15] , 
        \link_value_i[14] , \link_value_i[13] , \link_value_i[12] , 
        \link_value_i[11] , \link_value_i[10] , \link_value_i[9] , 
        \link_value_i[8] , \link_value_i[7] , \link_value_i[6] , 
        \link_value_i[5] , \link_value_i[4] , \link_value_i[3] , 
        \link_value_i[2] , \link_value_i[1] , \link_value_i[0] }) );
  mux21_NBIT32_0 jreg_mux21 ( .A(A_inALU_i), .B({\resAdd1_i[31] , 
        \resAdd1_i[30] , \resAdd1_i[29] , \resAdd1_i[28] , \resAdd1_i[27] , 
        \resAdd1_i[26] , \resAdd1_i[25] , \resAdd1_i[24] , \resAdd1_i[23] , 
        \resAdd1_i[22] , \resAdd1_i[21] , \resAdd1_i[20] , \resAdd1_i[19] , 
        \resAdd1_i[18] , \resAdd1_i[17] , \resAdd1_i[16] , \resAdd1_i[15] , 
        \resAdd1_i[14] , \resAdd1_i[13] , \resAdd1_i[12] , \resAdd1_i[11] , 
        \resAdd1_i[10] , \resAdd1_i[9] , \resAdd1_i[8] , \resAdd1_i[7] , 
        \resAdd1_i[6] , \resAdd1_i[5] , \resAdd1_i[4] , \resAdd1_i[3] , 
        \resAdd1_i[2] , \resAdd1_i[1] , \resAdd1_i[0] }), .S(controls_in_20), 
        .Y(toPC1) );
  mux21_NBIT32_5 link_mux21 ( .A({\link_value_i[31] , \link_value_i[30] , 
        \link_value_i[29] , \link_value_i[28] , \link_value_i[27] , 
        \link_value_i[26] , \link_value_i[25] , \link_value_i[24] , 
        \link_value_i[23] , \link_value_i[22] , \link_value_i[21] , 
        \link_value_i[20] , \link_value_i[19] , \link_value_i[18] , 
        \link_value_i[17] , \link_value_i[16] , \link_value_i[15] , 
        \link_value_i[14] , \link_value_i[13] , \link_value_i[12] , 
        \link_value_i[11] , \link_value_i[10] , \link_value_i[9] , 
        \link_value_i[8] , \link_value_i[7] , \link_value_i[6] , 
        \link_value_i[5] , \link_value_i[4] , \link_value_i[3] , 
        \link_value_i[2] , \link_value_i[1] , \link_value_i[0] }), .B(
        res_outALU_i), .S(\controls_in[18] ), .Y({\link2lhi_wire_i[31] , 
        \link2lhi_wire_i[30] , \link2lhi_wire_i[29] , \link2lhi_wire_i[28] , 
        \link2lhi_wire_i[27] , \link2lhi_wire_i[26] , \link2lhi_wire_i[25] , 
        \link2lhi_wire_i[24] , \link2lhi_wire_i[23] , \link2lhi_wire_i[22] , 
        \link2lhi_wire_i[21] , \link2lhi_wire_i[20] , \link2lhi_wire_i[19] , 
        \link2lhi_wire_i[18] , \link2lhi_wire_i[17] , \link2lhi_wire_i[16] , 
        \link2lhi_wire_i[15] , \link2lhi_wire_i[14] , \link2lhi_wire_i[13] , 
        \link2lhi_wire_i[12] , \link2lhi_wire_i[11] , \link2lhi_wire_i[10] , 
        \link2lhi_wire_i[9] , \link2lhi_wire_i[8] , \link2lhi_wire_i[7] , 
        \link2lhi_wire_i[6] , \link2lhi_wire_i[5] , \link2lhi_wire_i[4] , 
        \link2lhi_wire_i[3] , \link2lhi_wire_i[2] , \link2lhi_wire_i[1] , 
        \link2lhi_wire_i[0] }) );
  mux21_NBIT32_4 lhi_mux21 ( .A({lhi_value_i[31:16], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\link2lhi_wire_i[31] , \link2lhi_wire_i[30] , \link2lhi_wire_i[29] , 
        \link2lhi_wire_i[28] , \link2lhi_wire_i[27] , \link2lhi_wire_i[26] , 
        \link2lhi_wire_i[25] , \link2lhi_wire_i[24] , \link2lhi_wire_i[23] , 
        \link2lhi_wire_i[22] , \link2lhi_wire_i[21] , \link2lhi_wire_i[20] , 
        \link2lhi_wire_i[19] , \link2lhi_wire_i[18] , \link2lhi_wire_i[17] , 
        \link2lhi_wire_i[16] , \link2lhi_wire_i[15] , \link2lhi_wire_i[14] , 
        \link2lhi_wire_i[13] , \link2lhi_wire_i[12] , \link2lhi_wire_i[11] , 
        \link2lhi_wire_i[10] , \link2lhi_wire_i[9] , \link2lhi_wire_i[8] , 
        \link2lhi_wire_i[7] , \link2lhi_wire_i[6] , \link2lhi_wire_i[5] , 
        \link2lhi_wire_i[4] , \link2lhi_wire_i[3] , \link2lhi_wire_i[2] , 
        \link2lhi_wire_i[1] , \link2lhi_wire_i[0] }), .S(controls_in_17), .Y({
        \lhi2mov_wire_i[31] , \lhi2mov_wire_i[30] , \lhi2mov_wire_i[29] , 
        \lhi2mov_wire_i[28] , \lhi2mov_wire_i[27] , \lhi2mov_wire_i[26] , 
        \lhi2mov_wire_i[25] , \lhi2mov_wire_i[24] , \lhi2mov_wire_i[23] , 
        \lhi2mov_wire_i[22] , \lhi2mov_wire_i[21] , \lhi2mov_wire_i[20] , 
        \lhi2mov_wire_i[19] , \lhi2mov_wire_i[18] , \lhi2mov_wire_i[17] , 
        \lhi2mov_wire_i[16] , \lhi2mov_wire_i[15] , \lhi2mov_wire_i[14] , 
        \lhi2mov_wire_i[13] , \lhi2mov_wire_i[12] , \lhi2mov_wire_i[11] , 
        \lhi2mov_wire_i[10] , \lhi2mov_wire_i[9] , \lhi2mov_wire_i[8] , 
        \lhi2mov_wire_i[7] , \lhi2mov_wire_i[6] , \lhi2mov_wire_i[5] , 
        \lhi2mov_wire_i[4] , \lhi2mov_wire_i[3] , \lhi2mov_wire_i[2] , 
        \lhi2mov_wire_i[1] , \lhi2mov_wire_i[0] }) );
  mux21_NBIT5_0 regaddr_mux21 ( .A(rd_inst), .B(rt_inst), .S(controls_in_16), 
        .Y(addrRF) );
  mux21_NBIT32_3 movs2i_mux21 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        psw_status_i[1:0]}), .B({\lhi2mov_wire_i[31] , \lhi2mov_wire_i[30] , 
        \lhi2mov_wire_i[29] , \lhi2mov_wire_i[28] , \lhi2mov_wire_i[27] , 
        \lhi2mov_wire_i[26] , \lhi2mov_wire_i[25] , \lhi2mov_wire_i[24] , 
        \lhi2mov_wire_i[23] , \lhi2mov_wire_i[22] , \lhi2mov_wire_i[21] , 
        \lhi2mov_wire_i[20] , \lhi2mov_wire_i[19] , \lhi2mov_wire_i[18] , 
        \lhi2mov_wire_i[17] , \lhi2mov_wire_i[16] , \lhi2mov_wire_i[15] , 
        \lhi2mov_wire_i[14] , \lhi2mov_wire_i[13] , \lhi2mov_wire_i[12] , 
        \lhi2mov_wire_i[11] , \lhi2mov_wire_i[10] , \lhi2mov_wire_i[9] , 
        \lhi2mov_wire_i[8] , \lhi2mov_wire_i[7] , \lhi2mov_wire_i[6] , 
        \lhi2mov_wire_i[5] , \lhi2mov_wire_i[4] , \lhi2mov_wire_i[3] , 
        \lhi2mov_wire_i[2] , \lhi2mov_wire_i[1] , \lhi2mov_wire_i[0] }), .S(
        controls_in_15), .Y(addrMem) );
  mux21_NBIT32_2 alusrc_mux21 ( .A(ext15_0), .B(writeData), .S(controls_in_14), 
        .Y(B_inALU_i) );
  mux41_NBIT32_0 oprnd1_mux41 ( .a(op_A), .b(forw_dataWB), .c(forw_dataMEM), 
        .s(forwardA_i), .y(A_inALU_i) );
  mux41_NBIT32_1 oprnd2_mux41 ( .a(op_B), .b(forw_dataWB), .c(forw_dataMEM), 
        .s(forwardB_i), .y(writeData) );
  concat16 concatenate16 ( .string16(inst15_0), .string32({lhi_value_i[31:16], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15}) );
  forward forwarding_unit ( .rt_addr_IDEX(rt_inst), .rs_addr_IDEX(rs_inst), 
        .rd_addr_EXMEM(RFaddr_MEM), .rd_addr_MEMWB(RFaddr_WB), 
        .regwrite_EXMEM(regwriteMEM), .regwrite_MEMWB(regwriteWB), .forwardA(
        forwardA_i), .forwardB(forwardB_i) );
  branch_circ branch_circuit ( .branch_type(controls_in_19), .zero(zero_i), 
        .branch_taken(branchTaken) );
  PSWreg PSW ( .rst(rst), .clk(clk), .unaligned(unaligned), .ovf(ovf_i), 
        .status({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, psw_status_i[1:0]}) );
  ALU EXALU ( .alu_op(controls_in[4:0]), .a(A_inALU_i), .b(B_inALU_i), .ovf(
        ovf_i), .zero(zero_i), .res(res_outALU_i) );
endmodule


module idex_reg ( cw_to_ex_dec, jump_address_dec, pc_4_dec, read_data_1_dec, 
        read_data_2_dec, immediate_ext_dec, immediate_dec, rt_dec, rd_dec, 
        rs_dec, clk, rst, cw_to_ex, jump_address, pc_4, read_data_1, 
        read_data_2, immediate_ext, immediate, rt, rd, rs );
  input [21:0] cw_to_ex_dec;
  input [31:0] jump_address_dec;
  input [31:0] pc_4_dec;
  input [31:0] read_data_1_dec;
  input [31:0] read_data_2_dec;
  input [31:0] immediate_ext_dec;
  input [15:0] immediate_dec;
  input [4:0] rt_dec;
  input [4:0] rd_dec;
  input [4:0] rs_dec;
  output [21:0] cw_to_ex;
  output [31:0] jump_address;
  output [31:0] pc_4;
  output [31:0] read_data_1;
  output [31:0] read_data_2;
  output [31:0] immediate_ext;
  output [15:0] immediate;
  output [4:0] rt;
  output [4:0] rd;
  output [4:0] rs;
  input clk, rst;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, n215, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259;

  DFF_X1 \rs_reg[4]  ( .D(N215), .CK(clk), .Q(rs[4]) );
  DFF_X1 \rs_reg[3]  ( .D(N214), .CK(clk), .Q(rs[3]) );
  DFF_X1 \rs_reg[2]  ( .D(N213), .CK(clk), .Q(rs[2]) );
  DFF_X1 \rs_reg[1]  ( .D(N212), .CK(clk), .Q(rs[1]) );
  DFF_X1 \rs_reg[0]  ( .D(N211), .CK(clk), .Q(rs[0]) );
  DFF_X1 \cw_to_ex_reg[21]  ( .D(N24), .CK(clk), .Q(cw_to_ex[21]) );
  DFF_X1 \cw_to_ex_reg[20]  ( .D(N23), .CK(clk), .Q(cw_to_ex[20]) );
  DFF_X1 \cw_to_ex_reg[19]  ( .D(N22), .CK(clk), .Q(cw_to_ex[19]) );
  DFF_X1 \cw_to_ex_reg[18]  ( .D(N21), .CK(clk), .Q(cw_to_ex[18]) );
  DFF_X1 \cw_to_ex_reg[17]  ( .D(N20), .CK(clk), .Q(cw_to_ex[17]) );
  DFF_X1 \cw_to_ex_reg[16]  ( .D(N19), .CK(clk), .Q(cw_to_ex[16]) );
  DFF_X1 \cw_to_ex_reg[15]  ( .D(N18), .CK(clk), .Q(cw_to_ex[15]) );
  DFF_X1 \cw_to_ex_reg[14]  ( .D(N17), .CK(clk), .Q(cw_to_ex[14]) );
  DFF_X1 \cw_to_ex_reg[13]  ( .D(N16), .CK(clk), .Q(cw_to_ex[13]) );
  DFF_X1 \cw_to_ex_reg[12]  ( .D(N15), .CK(clk), .Q(cw_to_ex[12]) );
  DFF_X1 \cw_to_ex_reg[11]  ( .D(N14), .CK(clk), .Q(cw_to_ex[11]) );
  DFF_X1 \cw_to_ex_reg[10]  ( .D(N13), .CK(clk), .Q(cw_to_ex[10]) );
  DFF_X1 \cw_to_ex_reg[9]  ( .D(N12), .CK(clk), .Q(cw_to_ex[9]) );
  DFF_X1 \cw_to_ex_reg[8]  ( .D(N11), .CK(clk), .Q(cw_to_ex[8]) );
  DFF_X1 \cw_to_ex_reg[7]  ( .D(N10), .CK(clk), .Q(cw_to_ex[7]) );
  DFF_X1 \cw_to_ex_reg[6]  ( .D(N9), .CK(clk), .Q(cw_to_ex[6]) );
  DFF_X1 \cw_to_ex_reg[5]  ( .D(N8), .CK(clk), .Q(cw_to_ex[5]) );
  DFF_X1 \cw_to_ex_reg[4]  ( .D(N7), .CK(clk), .Q(cw_to_ex[4]) );
  DFF_X1 \cw_to_ex_reg[3]  ( .D(N6), .CK(clk), .Q(cw_to_ex[3]) );
  DFF_X1 \cw_to_ex_reg[2]  ( .D(N5), .CK(clk), .Q(cw_to_ex[2]) );
  DFF_X1 \cw_to_ex_reg[1]  ( .D(N4), .CK(clk), .Q(cw_to_ex[1]) );
  DFF_X1 \cw_to_ex_reg[0]  ( .D(N3), .CK(clk), .Q(cw_to_ex[0]) );
  DFF_X1 \jump_address_reg[31]  ( .D(N56), .CK(clk), .Q(jump_address[31]) );
  DFF_X1 \jump_address_reg[30]  ( .D(N55), .CK(clk), .Q(jump_address[30]) );
  DFF_X1 \jump_address_reg[29]  ( .D(N54), .CK(clk), .Q(jump_address[29]) );
  DFF_X1 \jump_address_reg[28]  ( .D(N53), .CK(clk), .Q(jump_address[28]) );
  DFF_X1 \jump_address_reg[27]  ( .D(N52), .CK(clk), .Q(jump_address[27]) );
  DFF_X1 \jump_address_reg[26]  ( .D(N51), .CK(clk), .Q(jump_address[26]) );
  DFF_X1 \jump_address_reg[25]  ( .D(N50), .CK(clk), .Q(jump_address[25]) );
  DFF_X1 \jump_address_reg[24]  ( .D(N49), .CK(clk), .Q(jump_address[24]) );
  DFF_X1 \jump_address_reg[23]  ( .D(N48), .CK(clk), .Q(jump_address[23]) );
  DFF_X1 \jump_address_reg[22]  ( .D(N47), .CK(clk), .Q(jump_address[22]) );
  DFF_X1 \jump_address_reg[21]  ( .D(N46), .CK(clk), .Q(jump_address[21]) );
  DFF_X1 \jump_address_reg[20]  ( .D(N45), .CK(clk), .Q(jump_address[20]) );
  DFF_X1 \jump_address_reg[19]  ( .D(N44), .CK(clk), .Q(jump_address[19]) );
  DFF_X1 \jump_address_reg[18]  ( .D(N43), .CK(clk), .Q(jump_address[18]) );
  DFF_X1 \jump_address_reg[17]  ( .D(N42), .CK(clk), .Q(jump_address[17]) );
  DFF_X1 \jump_address_reg[16]  ( .D(N41), .CK(clk), .Q(jump_address[16]) );
  DFF_X1 \jump_address_reg[15]  ( .D(N40), .CK(clk), .Q(jump_address[15]) );
  DFF_X1 \jump_address_reg[14]  ( .D(N39), .CK(clk), .Q(jump_address[14]) );
  DFF_X1 \jump_address_reg[13]  ( .D(N38), .CK(clk), .Q(jump_address[13]) );
  DFF_X1 \jump_address_reg[12]  ( .D(N37), .CK(clk), .Q(jump_address[12]) );
  DFF_X1 \jump_address_reg[11]  ( .D(N36), .CK(clk), .Q(jump_address[11]) );
  DFF_X1 \jump_address_reg[10]  ( .D(N35), .CK(clk), .Q(jump_address[10]) );
  DFF_X1 \jump_address_reg[9]  ( .D(N34), .CK(clk), .Q(jump_address[9]) );
  DFF_X1 \jump_address_reg[8]  ( .D(N33), .CK(clk), .Q(jump_address[8]) );
  DFF_X1 \jump_address_reg[7]  ( .D(N32), .CK(clk), .Q(jump_address[7]) );
  DFF_X1 \jump_address_reg[6]  ( .D(N31), .CK(clk), .Q(jump_address[6]) );
  DFF_X1 \jump_address_reg[5]  ( .D(N30), .CK(clk), .Q(jump_address[5]) );
  DFF_X1 \jump_address_reg[4]  ( .D(N29), .CK(clk), .Q(jump_address[4]) );
  DFF_X1 \jump_address_reg[3]  ( .D(N28), .CK(clk), .Q(jump_address[3]) );
  DFF_X1 \jump_address_reg[2]  ( .D(N27), .CK(clk), .Q(jump_address[2]) );
  DFF_X1 \jump_address_reg[1]  ( .D(N26), .CK(clk), .Q(jump_address[1]) );
  DFF_X1 \jump_address_reg[0]  ( .D(N25), .CK(clk), .Q(jump_address[0]) );
  DFF_X1 \pc_4_reg[31]  ( .D(N88), .CK(clk), .Q(pc_4[31]) );
  DFF_X1 \pc_4_reg[30]  ( .D(N87), .CK(clk), .Q(pc_4[30]) );
  DFF_X1 \pc_4_reg[29]  ( .D(N86), .CK(clk), .Q(pc_4[29]) );
  DFF_X1 \pc_4_reg[28]  ( .D(N85), .CK(clk), .Q(pc_4[28]) );
  DFF_X1 \pc_4_reg[27]  ( .D(N84), .CK(clk), .Q(pc_4[27]) );
  DFF_X1 \pc_4_reg[26]  ( .D(N83), .CK(clk), .Q(pc_4[26]) );
  DFF_X1 \pc_4_reg[25]  ( .D(N82), .CK(clk), .Q(pc_4[25]) );
  DFF_X1 \pc_4_reg[24]  ( .D(N81), .CK(clk), .Q(pc_4[24]) );
  DFF_X1 \pc_4_reg[23]  ( .D(N80), .CK(clk), .Q(pc_4[23]) );
  DFF_X1 \pc_4_reg[22]  ( .D(N79), .CK(clk), .Q(pc_4[22]) );
  DFF_X1 \pc_4_reg[21]  ( .D(N78), .CK(clk), .Q(pc_4[21]) );
  DFF_X1 \pc_4_reg[20]  ( .D(N77), .CK(clk), .Q(pc_4[20]) );
  DFF_X1 \pc_4_reg[19]  ( .D(N76), .CK(clk), .Q(pc_4[19]) );
  DFF_X1 \pc_4_reg[18]  ( .D(N75), .CK(clk), .Q(pc_4[18]) );
  DFF_X1 \pc_4_reg[17]  ( .D(N74), .CK(clk), .Q(pc_4[17]) );
  DFF_X1 \pc_4_reg[16]  ( .D(N73), .CK(clk), .Q(pc_4[16]) );
  DFF_X1 \pc_4_reg[15]  ( .D(N72), .CK(clk), .Q(pc_4[15]) );
  DFF_X1 \pc_4_reg[14]  ( .D(N71), .CK(clk), .Q(pc_4[14]) );
  DFF_X1 \pc_4_reg[13]  ( .D(N70), .CK(clk), .Q(pc_4[13]) );
  DFF_X1 \pc_4_reg[12]  ( .D(N69), .CK(clk), .Q(pc_4[12]) );
  DFF_X1 \pc_4_reg[11]  ( .D(N68), .CK(clk), .Q(pc_4[11]) );
  DFF_X1 \pc_4_reg[10]  ( .D(N67), .CK(clk), .Q(pc_4[10]) );
  DFF_X1 \pc_4_reg[9]  ( .D(N66), .CK(clk), .Q(pc_4[9]) );
  DFF_X1 \pc_4_reg[8]  ( .D(N65), .CK(clk), .Q(pc_4[8]) );
  DFF_X1 \pc_4_reg[7]  ( .D(N64), .CK(clk), .Q(pc_4[7]) );
  DFF_X1 \pc_4_reg[6]  ( .D(N63), .CK(clk), .Q(pc_4[6]) );
  DFF_X1 \pc_4_reg[5]  ( .D(N62), .CK(clk), .Q(pc_4[5]) );
  DFF_X1 \pc_4_reg[4]  ( .D(N61), .CK(clk), .Q(pc_4[4]) );
  DFF_X1 \pc_4_reg[3]  ( .D(N60), .CK(clk), .Q(pc_4[3]) );
  DFF_X1 \pc_4_reg[2]  ( .D(N59), .CK(clk), .Q(pc_4[2]) );
  DFF_X1 \pc_4_reg[1]  ( .D(N58), .CK(clk), .Q(pc_4[1]) );
  DFF_X1 \pc_4_reg[0]  ( .D(N57), .CK(clk), .Q(pc_4[0]) );
  DFF_X1 \read_data_1_reg[31]  ( .D(N120), .CK(clk), .Q(read_data_1[31]) );
  DFF_X1 \read_data_1_reg[30]  ( .D(N119), .CK(clk), .Q(read_data_1[30]) );
  DFF_X1 \read_data_1_reg[29]  ( .D(N118), .CK(clk), .Q(read_data_1[29]) );
  DFF_X1 \read_data_1_reg[28]  ( .D(N117), .CK(clk), .Q(read_data_1[28]) );
  DFF_X1 \read_data_1_reg[27]  ( .D(N116), .CK(clk), .Q(read_data_1[27]) );
  DFF_X1 \read_data_1_reg[26]  ( .D(N115), .CK(clk), .Q(read_data_1[26]) );
  DFF_X1 \read_data_1_reg[25]  ( .D(N114), .CK(clk), .Q(read_data_1[25]) );
  DFF_X1 \read_data_1_reg[24]  ( .D(N113), .CK(clk), .Q(read_data_1[24]) );
  DFF_X1 \read_data_1_reg[23]  ( .D(N112), .CK(clk), .Q(read_data_1[23]) );
  DFF_X1 \read_data_1_reg[22]  ( .D(N111), .CK(clk), .Q(read_data_1[22]) );
  DFF_X1 \read_data_1_reg[21]  ( .D(N110), .CK(clk), .Q(read_data_1[21]) );
  DFF_X1 \read_data_1_reg[20]  ( .D(N109), .CK(clk), .Q(read_data_1[20]) );
  DFF_X1 \read_data_1_reg[19]  ( .D(N108), .CK(clk), .Q(read_data_1[19]) );
  DFF_X1 \read_data_1_reg[18]  ( .D(N107), .CK(clk), .Q(read_data_1[18]) );
  DFF_X1 \read_data_1_reg[17]  ( .D(N106), .CK(clk), .Q(read_data_1[17]) );
  DFF_X1 \read_data_1_reg[16]  ( .D(N105), .CK(clk), .Q(read_data_1[16]) );
  DFF_X1 \read_data_1_reg[15]  ( .D(N104), .CK(clk), .Q(read_data_1[15]) );
  DFF_X1 \read_data_1_reg[14]  ( .D(N103), .CK(clk), .Q(read_data_1[14]) );
  DFF_X1 \read_data_1_reg[13]  ( .D(N102), .CK(clk), .Q(read_data_1[13]) );
  DFF_X1 \read_data_1_reg[12]  ( .D(N101), .CK(clk), .Q(read_data_1[12]) );
  DFF_X1 \read_data_1_reg[11]  ( .D(N100), .CK(clk), .Q(read_data_1[11]) );
  DFF_X1 \read_data_1_reg[10]  ( .D(N99), .CK(clk), .Q(read_data_1[10]) );
  DFF_X1 \read_data_1_reg[9]  ( .D(N98), .CK(clk), .Q(read_data_1[9]) );
  DFF_X1 \read_data_1_reg[8]  ( .D(N97), .CK(clk), .Q(read_data_1[8]) );
  DFF_X1 \read_data_1_reg[7]  ( .D(N96), .CK(clk), .Q(read_data_1[7]) );
  DFF_X1 \read_data_1_reg[6]  ( .D(N95), .CK(clk), .Q(read_data_1[6]) );
  DFF_X1 \read_data_1_reg[5]  ( .D(N94), .CK(clk), .Q(read_data_1[5]) );
  DFF_X1 \read_data_1_reg[4]  ( .D(N93), .CK(clk), .Q(read_data_1[4]) );
  DFF_X1 \read_data_1_reg[3]  ( .D(N92), .CK(clk), .Q(read_data_1[3]) );
  DFF_X1 \read_data_1_reg[2]  ( .D(N91), .CK(clk), .Q(read_data_1[2]) );
  DFF_X1 \read_data_1_reg[1]  ( .D(N90), .CK(clk), .Q(read_data_1[1]) );
  DFF_X1 \read_data_1_reg[0]  ( .D(N89), .CK(clk), .Q(read_data_1[0]) );
  DFF_X1 \read_data_2_reg[31]  ( .D(N152), .CK(clk), .Q(read_data_2[31]) );
  DFF_X1 \read_data_2_reg[30]  ( .D(N151), .CK(clk), .Q(read_data_2[30]) );
  DFF_X1 \read_data_2_reg[29]  ( .D(N150), .CK(clk), .Q(read_data_2[29]) );
  DFF_X1 \read_data_2_reg[28]  ( .D(N149), .CK(clk), .Q(read_data_2[28]) );
  DFF_X1 \read_data_2_reg[27]  ( .D(N148), .CK(clk), .Q(read_data_2[27]) );
  DFF_X1 \read_data_2_reg[26]  ( .D(N147), .CK(clk), .Q(read_data_2[26]) );
  DFF_X1 \read_data_2_reg[25]  ( .D(N146), .CK(clk), .Q(read_data_2[25]) );
  DFF_X1 \read_data_2_reg[24]  ( .D(N145), .CK(clk), .Q(read_data_2[24]) );
  DFF_X1 \read_data_2_reg[23]  ( .D(N144), .CK(clk), .Q(read_data_2[23]) );
  DFF_X1 \read_data_2_reg[22]  ( .D(N143), .CK(clk), .Q(read_data_2[22]) );
  DFF_X1 \read_data_2_reg[21]  ( .D(N142), .CK(clk), .Q(read_data_2[21]) );
  DFF_X1 \read_data_2_reg[20]  ( .D(N141), .CK(clk), .Q(read_data_2[20]) );
  DFF_X1 \read_data_2_reg[19]  ( .D(N140), .CK(clk), .Q(read_data_2[19]) );
  DFF_X1 \read_data_2_reg[18]  ( .D(N139), .CK(clk), .Q(read_data_2[18]) );
  DFF_X1 \read_data_2_reg[17]  ( .D(N138), .CK(clk), .Q(read_data_2[17]) );
  DFF_X1 \read_data_2_reg[16]  ( .D(N137), .CK(clk), .Q(read_data_2[16]) );
  DFF_X1 \read_data_2_reg[15]  ( .D(N136), .CK(clk), .Q(read_data_2[15]) );
  DFF_X1 \read_data_2_reg[14]  ( .D(N135), .CK(clk), .Q(read_data_2[14]) );
  DFF_X1 \read_data_2_reg[13]  ( .D(N134), .CK(clk), .Q(read_data_2[13]) );
  DFF_X1 \read_data_2_reg[12]  ( .D(N133), .CK(clk), .Q(read_data_2[12]) );
  DFF_X1 \read_data_2_reg[11]  ( .D(N132), .CK(clk), .Q(read_data_2[11]) );
  DFF_X1 \read_data_2_reg[10]  ( .D(N131), .CK(clk), .Q(read_data_2[10]) );
  DFF_X1 \read_data_2_reg[9]  ( .D(N130), .CK(clk), .Q(read_data_2[9]) );
  DFF_X1 \read_data_2_reg[8]  ( .D(N129), .CK(clk), .Q(read_data_2[8]) );
  DFF_X1 \read_data_2_reg[7]  ( .D(N128), .CK(clk), .Q(read_data_2[7]) );
  DFF_X1 \read_data_2_reg[6]  ( .D(N127), .CK(clk), .Q(read_data_2[6]) );
  DFF_X1 \read_data_2_reg[5]  ( .D(N126), .CK(clk), .Q(read_data_2[5]) );
  DFF_X1 \read_data_2_reg[4]  ( .D(N125), .CK(clk), .Q(read_data_2[4]) );
  DFF_X1 \read_data_2_reg[3]  ( .D(N124), .CK(clk), .Q(read_data_2[3]) );
  DFF_X1 \read_data_2_reg[2]  ( .D(N123), .CK(clk), .Q(read_data_2[2]) );
  DFF_X1 \read_data_2_reg[1]  ( .D(N122), .CK(clk), .Q(read_data_2[1]) );
  DFF_X1 \read_data_2_reg[0]  ( .D(N121), .CK(clk), .Q(read_data_2[0]) );
  DFF_X1 \immediate_ext_reg[31]  ( .D(N184), .CK(clk), .Q(immediate_ext[31])
         );
  DFF_X1 \immediate_ext_reg[30]  ( .D(N183), .CK(clk), .Q(immediate_ext[30])
         );
  DFF_X1 \immediate_ext_reg[29]  ( .D(N182), .CK(clk), .Q(immediate_ext[29])
         );
  DFF_X1 \immediate_ext_reg[28]  ( .D(N181), .CK(clk), .Q(immediate_ext[28])
         );
  DFF_X1 \immediate_ext_reg[27]  ( .D(N180), .CK(clk), .Q(immediate_ext[27])
         );
  DFF_X1 \immediate_ext_reg[26]  ( .D(N179), .CK(clk), .Q(immediate_ext[26])
         );
  DFF_X1 \immediate_ext_reg[25]  ( .D(N178), .CK(clk), .Q(immediate_ext[25])
         );
  DFF_X1 \immediate_ext_reg[24]  ( .D(N177), .CK(clk), .Q(immediate_ext[24])
         );
  DFF_X1 \immediate_ext_reg[23]  ( .D(N176), .CK(clk), .Q(immediate_ext[23])
         );
  DFF_X1 \immediate_ext_reg[22]  ( .D(N175), .CK(clk), .Q(immediate_ext[22])
         );
  DFF_X1 \immediate_ext_reg[21]  ( .D(N174), .CK(clk), .Q(immediate_ext[21])
         );
  DFF_X1 \immediate_ext_reg[20]  ( .D(N173), .CK(clk), .Q(immediate_ext[20])
         );
  DFF_X1 \immediate_ext_reg[19]  ( .D(N172), .CK(clk), .Q(immediate_ext[19])
         );
  DFF_X1 \immediate_ext_reg[18]  ( .D(N171), .CK(clk), .Q(immediate_ext[18])
         );
  DFF_X1 \immediate_ext_reg[17]  ( .D(N170), .CK(clk), .Q(immediate_ext[17])
         );
  DFF_X1 \immediate_ext_reg[16]  ( .D(N169), .CK(clk), .Q(immediate_ext[16])
         );
  DFF_X1 \immediate_ext_reg[15]  ( .D(N168), .CK(clk), .Q(immediate_ext[15])
         );
  DFF_X1 \immediate_ext_reg[14]  ( .D(N167), .CK(clk), .Q(immediate_ext[14])
         );
  DFF_X1 \immediate_ext_reg[13]  ( .D(N166), .CK(clk), .Q(immediate_ext[13])
         );
  DFF_X1 \immediate_ext_reg[12]  ( .D(N165), .CK(clk), .Q(immediate_ext[12])
         );
  DFF_X1 \immediate_ext_reg[11]  ( .D(N164), .CK(clk), .Q(immediate_ext[11])
         );
  DFF_X1 \immediate_ext_reg[10]  ( .D(N163), .CK(clk), .Q(immediate_ext[10])
         );
  DFF_X1 \immediate_ext_reg[9]  ( .D(N162), .CK(clk), .Q(immediate_ext[9]) );
  DFF_X1 \immediate_ext_reg[8]  ( .D(N161), .CK(clk), .Q(immediate_ext[8]) );
  DFF_X1 \immediate_ext_reg[7]  ( .D(N160), .CK(clk), .Q(immediate_ext[7]) );
  DFF_X1 \immediate_ext_reg[6]  ( .D(N159), .CK(clk), .Q(immediate_ext[6]) );
  DFF_X1 \immediate_ext_reg[5]  ( .D(N158), .CK(clk), .Q(immediate_ext[5]) );
  DFF_X1 \immediate_ext_reg[4]  ( .D(N157), .CK(clk), .Q(immediate_ext[4]) );
  DFF_X1 \immediate_ext_reg[3]  ( .D(N156), .CK(clk), .Q(immediate_ext[3]) );
  DFF_X1 \immediate_ext_reg[2]  ( .D(N155), .CK(clk), .Q(immediate_ext[2]) );
  DFF_X1 \immediate_ext_reg[1]  ( .D(N154), .CK(clk), .Q(immediate_ext[1]) );
  DFF_X1 \immediate_ext_reg[0]  ( .D(N153), .CK(clk), .Q(immediate_ext[0]) );
  DFF_X1 \immediate_reg[15]  ( .D(N200), .CK(clk), .Q(immediate[15]) );
  DFF_X1 \immediate_reg[14]  ( .D(N199), .CK(clk), .Q(immediate[14]) );
  DFF_X1 \immediate_reg[13]  ( .D(N198), .CK(clk), .Q(immediate[13]) );
  DFF_X1 \immediate_reg[12]  ( .D(N197), .CK(clk), .Q(immediate[12]) );
  DFF_X1 \immediate_reg[11]  ( .D(N196), .CK(clk), .Q(immediate[11]) );
  DFF_X1 \immediate_reg[10]  ( .D(N195), .CK(clk), .Q(immediate[10]) );
  DFF_X1 \immediate_reg[9]  ( .D(N194), .CK(clk), .Q(immediate[9]) );
  DFF_X1 \immediate_reg[8]  ( .D(N193), .CK(clk), .Q(immediate[8]) );
  DFF_X1 \immediate_reg[7]  ( .D(N192), .CK(clk), .Q(immediate[7]) );
  DFF_X1 \immediate_reg[6]  ( .D(N191), .CK(clk), .Q(immediate[6]) );
  DFF_X1 \immediate_reg[5]  ( .D(N190), .CK(clk), .Q(immediate[5]) );
  DFF_X1 \immediate_reg[4]  ( .D(N189), .CK(clk), .Q(immediate[4]) );
  DFF_X1 \immediate_reg[3]  ( .D(N188), .CK(clk), .Q(immediate[3]) );
  DFF_X1 \immediate_reg[2]  ( .D(N187), .CK(clk), .Q(immediate[2]) );
  DFF_X1 \immediate_reg[1]  ( .D(N186), .CK(clk), .Q(immediate[1]) );
  DFF_X1 \immediate_reg[0]  ( .D(N185), .CK(clk), .Q(immediate[0]) );
  DFF_X1 \rt_reg[4]  ( .D(N205), .CK(clk), .Q(rt[4]) );
  DFF_X1 \rt_reg[3]  ( .D(N204), .CK(clk), .Q(rt[3]) );
  DFF_X1 \rt_reg[2]  ( .D(N203), .CK(clk), .Q(rt[2]) );
  DFF_X1 \rt_reg[1]  ( .D(N202), .CK(clk), .Q(rt[1]) );
  DFF_X1 \rt_reg[0]  ( .D(N201), .CK(clk), .Q(rt[0]) );
  DFF_X1 \rd_reg[4]  ( .D(N210), .CK(clk), .Q(rd[4]) );
  DFF_X1 \rd_reg[3]  ( .D(N209), .CK(clk), .Q(rd[3]) );
  DFF_X1 \rd_reg[2]  ( .D(N208), .CK(clk), .Q(rd[2]) );
  DFF_X1 \rd_reg[1]  ( .D(N207), .CK(clk), .Q(rd[1]) );
  DFF_X1 \rd_reg[0]  ( .D(N206), .CK(clk), .Q(rd[0]) );
  BUF_X1 U3 ( .A(n240), .Z(n253) );
  BUF_X1 U4 ( .A(n241), .Z(n254) );
  BUF_X1 U5 ( .A(n241), .Z(n255) );
  BUF_X1 U6 ( .A(n241), .Z(n256) );
  BUF_X1 U7 ( .A(n241), .Z(n257) );
  BUF_X1 U8 ( .A(n241), .Z(n258) );
  BUF_X1 U9 ( .A(n239), .Z(n242) );
  BUF_X1 U10 ( .A(n239), .Z(n243) );
  BUF_X1 U11 ( .A(n239), .Z(n244) );
  BUF_X1 U12 ( .A(n239), .Z(n245) );
  BUF_X1 U13 ( .A(n239), .Z(n246) );
  BUF_X1 U14 ( .A(n239), .Z(n247) );
  BUF_X1 U15 ( .A(n240), .Z(n248) );
  BUF_X1 U16 ( .A(n240), .Z(n249) );
  BUF_X1 U17 ( .A(n240), .Z(n250) );
  BUF_X1 U18 ( .A(n240), .Z(n251) );
  BUF_X1 U19 ( .A(n240), .Z(n252) );
  BUF_X1 U20 ( .A(n241), .Z(n259) );
  AND2_X1 U21 ( .A1(cw_to_ex_dec[7]), .A2(n242), .ZN(N10) );
  AND2_X1 U22 ( .A1(cw_to_ex_dec[12]), .A2(n246), .ZN(N15) );
  AND2_X1 U23 ( .A1(cw_to_ex_dec[16]), .A2(n250), .ZN(N19) );
  AND2_X1 U24 ( .A1(cw_to_ex_dec[18]), .A2(n252), .ZN(N21) );
  AND2_X1 U25 ( .A1(read_data_2_dec[3]), .A2(n244), .ZN(N124) );
  AND2_X1 U26 ( .A1(read_data_2_dec[4]), .A2(n244), .ZN(N125) );
  AND2_X1 U27 ( .A1(read_data_2_dec[5]), .A2(n244), .ZN(N126) );
  AND2_X1 U28 ( .A1(read_data_2_dec[6]), .A2(n244), .ZN(N127) );
  AND2_X1 U29 ( .A1(read_data_2_dec[7]), .A2(n244), .ZN(N128) );
  AND2_X1 U30 ( .A1(read_data_2_dec[8]), .A2(n244), .ZN(N129) );
  AND2_X1 U31 ( .A1(read_data_2_dec[9]), .A2(n244), .ZN(N130) );
  AND2_X1 U32 ( .A1(read_data_2_dec[31]), .A2(n246), .ZN(N152) );
  AND2_X1 U33 ( .A1(read_data_2_dec[0]), .A2(n244), .ZN(N121) );
  AND2_X1 U34 ( .A1(read_data_2_dec[1]), .A2(n244), .ZN(N122) );
  AND2_X1 U35 ( .A1(read_data_2_dec[2]), .A2(n244), .ZN(N123) );
  AND2_X1 U36 ( .A1(read_data_2_dec[10]), .A2(n244), .ZN(N131) );
  AND2_X1 U37 ( .A1(read_data_2_dec[11]), .A2(n245), .ZN(N132) );
  AND2_X1 U38 ( .A1(read_data_2_dec[12]), .A2(n245), .ZN(N133) );
  AND2_X1 U39 ( .A1(read_data_2_dec[13]), .A2(n245), .ZN(N134) );
  AND2_X1 U40 ( .A1(read_data_2_dec[14]), .A2(n245), .ZN(N135) );
  AND2_X1 U41 ( .A1(read_data_2_dec[15]), .A2(n245), .ZN(N136) );
  AND2_X1 U42 ( .A1(read_data_2_dec[16]), .A2(n245), .ZN(N137) );
  AND2_X1 U43 ( .A1(read_data_2_dec[17]), .A2(n245), .ZN(N138) );
  AND2_X1 U44 ( .A1(read_data_2_dec[18]), .A2(n245), .ZN(N139) );
  AND2_X1 U45 ( .A1(read_data_2_dec[19]), .A2(n245), .ZN(N140) );
  AND2_X1 U46 ( .A1(read_data_2_dec[20]), .A2(n245), .ZN(N141) );
  AND2_X1 U47 ( .A1(read_data_2_dec[21]), .A2(n245), .ZN(N142) );
  AND2_X1 U48 ( .A1(read_data_2_dec[22]), .A2(n246), .ZN(N143) );
  AND2_X1 U49 ( .A1(read_data_2_dec[23]), .A2(n246), .ZN(N144) );
  AND2_X1 U50 ( .A1(read_data_2_dec[24]), .A2(n246), .ZN(N145) );
  AND2_X1 U51 ( .A1(read_data_2_dec[25]), .A2(n246), .ZN(N146) );
  AND2_X1 U52 ( .A1(read_data_2_dec[26]), .A2(n246), .ZN(N147) );
  AND2_X1 U53 ( .A1(read_data_2_dec[27]), .A2(n246), .ZN(N148) );
  AND2_X1 U54 ( .A1(read_data_2_dec[28]), .A2(n246), .ZN(N149) );
  AND2_X1 U55 ( .A1(read_data_2_dec[29]), .A2(n246), .ZN(N150) );
  AND2_X1 U56 ( .A1(read_data_2_dec[30]), .A2(n246), .ZN(N151) );
  BUF_X1 U57 ( .A(n215), .Z(n241) );
  BUF_X1 U58 ( .A(n215), .Z(n239) );
  BUF_X1 U59 ( .A(n215), .Z(n240) );
  AND2_X1 U60 ( .A1(immediate_ext_dec[16]), .A2(n248), .ZN(N169) );
  AND2_X1 U61 ( .A1(immediate_ext_dec[17]), .A2(n248), .ZN(N170) );
  AND2_X1 U62 ( .A1(immediate_ext_dec[18]), .A2(n248), .ZN(N171) );
  AND2_X1 U63 ( .A1(immediate_ext_dec[19]), .A2(n248), .ZN(N172) );
  AND2_X1 U64 ( .A1(immediate_ext_dec[20]), .A2(n248), .ZN(N173) );
  AND2_X1 U65 ( .A1(immediate_ext_dec[21]), .A2(n248), .ZN(N174) );
  AND2_X1 U66 ( .A1(immediate_ext_dec[22]), .A2(n248), .ZN(N175) );
  AND2_X1 U67 ( .A1(immediate_ext_dec[23]), .A2(n249), .ZN(N176) );
  AND2_X1 U68 ( .A1(immediate_ext_dec[24]), .A2(n249), .ZN(N177) );
  AND2_X1 U69 ( .A1(immediate_ext_dec[25]), .A2(n249), .ZN(N178) );
  AND2_X1 U70 ( .A1(immediate_ext_dec[26]), .A2(n249), .ZN(N179) );
  AND2_X1 U71 ( .A1(immediate_ext_dec[27]), .A2(n249), .ZN(N180) );
  AND2_X1 U72 ( .A1(immediate_ext_dec[28]), .A2(n249), .ZN(N181) );
  AND2_X1 U73 ( .A1(immediate_ext_dec[29]), .A2(n249), .ZN(N182) );
  AND2_X1 U74 ( .A1(immediate_ext_dec[30]), .A2(n249), .ZN(N183) );
  AND2_X1 U75 ( .A1(immediate_ext_dec[31]), .A2(n249), .ZN(N184) );
  AND2_X1 U76 ( .A1(cw_to_ex_dec[0]), .A2(n253), .ZN(N3) );
  AND2_X1 U77 ( .A1(cw_to_ex_dec[1]), .A2(n254), .ZN(N4) );
  AND2_X1 U78 ( .A1(cw_to_ex_dec[5]), .A2(n257), .ZN(N8) );
  AND2_X1 U79 ( .A1(cw_to_ex_dec[6]), .A2(n258), .ZN(N9) );
  AND2_X1 U80 ( .A1(cw_to_ex_dec[8]), .A2(n242), .ZN(N11) );
  AND2_X1 U81 ( .A1(cw_to_ex_dec[9]), .A2(n243), .ZN(N12) );
  AND2_X1 U82 ( .A1(cw_to_ex_dec[10]), .A2(n244), .ZN(N13) );
  AND2_X1 U83 ( .A1(cw_to_ex_dec[13]), .A2(n247), .ZN(N16) );
  AND2_X1 U84 ( .A1(cw_to_ex_dec[17]), .A2(n251), .ZN(N20) );
  AND2_X1 U85 ( .A1(cw_to_ex_dec[20]), .A2(n252), .ZN(N23) );
  AND2_X1 U86 ( .A1(cw_to_ex_dec[21]), .A2(n252), .ZN(N24) );
  AND2_X1 U87 ( .A1(immediate_dec[2]), .A2(n250), .ZN(N187) );
  AND2_X1 U88 ( .A1(immediate_ext_dec[2]), .A2(n247), .ZN(N155) );
  AND2_X1 U89 ( .A1(jump_address_dec[2]), .A2(n253), .ZN(N27) );
  INV_X1 U90 ( .A(rst), .ZN(n215) );
  AND2_X1 U91 ( .A1(jump_address_dec[25]), .A2(n255), .ZN(N50) );
  AND2_X1 U92 ( .A1(jump_address_dec[26]), .A2(n255), .ZN(N51) );
  AND2_X1 U93 ( .A1(jump_address_dec[27]), .A2(n255), .ZN(N52) );
  AND2_X1 U94 ( .A1(jump_address_dec[28]), .A2(n255), .ZN(N53) );
  AND2_X1 U95 ( .A1(jump_address_dec[29]), .A2(n255), .ZN(N54) );
  AND2_X1 U96 ( .A1(jump_address_dec[30]), .A2(n255), .ZN(N55) );
  AND2_X1 U97 ( .A1(jump_address_dec[31]), .A2(n255), .ZN(N56) );
  AND2_X1 U98 ( .A1(rs_dec[4]), .A2(n252), .ZN(N215) );
  AND2_X1 U99 ( .A1(rt_dec[2]), .A2(n251), .ZN(N203) );
  AND2_X1 U100 ( .A1(jump_address_dec[18]), .A2(n254), .ZN(N43) );
  AND2_X1 U101 ( .A1(immediate_dec[3]), .A2(n250), .ZN(N188) );
  AND2_X1 U102 ( .A1(immediate_ext_dec[3]), .A2(n247), .ZN(N156) );
  AND2_X1 U103 ( .A1(jump_address_dec[3]), .A2(n253), .ZN(N28) );
  AND2_X1 U104 ( .A1(immediate_dec[0]), .A2(n249), .ZN(N185) );
  AND2_X1 U105 ( .A1(immediate_ext_dec[0]), .A2(n246), .ZN(N153) );
  AND2_X1 U106 ( .A1(jump_address_dec[0]), .A2(n252), .ZN(N25) );
  AND2_X1 U107 ( .A1(jump_address_dec[23]), .A2(n255), .ZN(N48) );
  AND2_X1 U108 ( .A1(rs_dec[2]), .A2(n252), .ZN(N213) );
  AND2_X1 U109 ( .A1(immediate_dec[1]), .A2(n249), .ZN(N186) );
  AND2_X1 U110 ( .A1(immediate_ext_dec[1]), .A2(n247), .ZN(N154) );
  AND2_X1 U111 ( .A1(jump_address_dec[1]), .A2(n253), .ZN(N26) );
  AND2_X1 U112 ( .A1(immediate_dec[5]), .A2(n250), .ZN(N190) );
  AND2_X1 U113 ( .A1(immediate_ext_dec[5]), .A2(n247), .ZN(N158) );
  AND2_X1 U114 ( .A1(jump_address_dec[5]), .A2(n253), .ZN(N30) );
  AND2_X1 U115 ( .A1(jump_address_dec[22]), .A2(n254), .ZN(N47) );
  AND2_X1 U116 ( .A1(rs_dec[1]), .A2(n252), .ZN(N212) );
  AND2_X1 U117 ( .A1(rt_dec[4]), .A2(n251), .ZN(N205) );
  AND2_X1 U118 ( .A1(jump_address_dec[20]), .A2(n254), .ZN(N45) );
  AND2_X1 U119 ( .A1(rt_dec[1]), .A2(n251), .ZN(N202) );
  AND2_X1 U120 ( .A1(rt_dec[3]), .A2(n251), .ZN(N204) );
  AND2_X1 U121 ( .A1(jump_address_dec[17]), .A2(n254), .ZN(N42) );
  AND2_X1 U122 ( .A1(jump_address_dec[19]), .A2(n254), .ZN(N44) );
  AND2_X1 U123 ( .A1(jump_address_dec[21]), .A2(n254), .ZN(N46) );
  AND2_X1 U124 ( .A1(rs_dec[0]), .A2(n252), .ZN(N211) );
  AND2_X1 U125 ( .A1(jump_address_dec[24]), .A2(n255), .ZN(N49) );
  AND2_X1 U126 ( .A1(rs_dec[3]), .A2(n252), .ZN(N214) );
  AND2_X1 U127 ( .A1(immediate_dec[4]), .A2(n250), .ZN(N189) );
  AND2_X1 U128 ( .A1(immediate_ext_dec[4]), .A2(n247), .ZN(N157) );
  AND2_X1 U129 ( .A1(jump_address_dec[4]), .A2(n253), .ZN(N29) );
  AND2_X1 U130 ( .A1(rt_dec[0]), .A2(n251), .ZN(N201) );
  AND2_X1 U131 ( .A1(jump_address_dec[16]), .A2(n254), .ZN(N41) );
  AND2_X1 U132 ( .A1(rd_dec[4]), .A2(n252), .ZN(N210) );
  AND2_X1 U133 ( .A1(immediate_dec[15]), .A2(n251), .ZN(N200) );
  AND2_X1 U134 ( .A1(immediate_ext_dec[15]), .A2(n248), .ZN(N168) );
  AND2_X1 U135 ( .A1(jump_address_dec[15]), .A2(n254), .ZN(N40) );
  AND2_X1 U136 ( .A1(immediate_dec[6]), .A2(n250), .ZN(N191) );
  AND2_X1 U137 ( .A1(immediate_ext_dec[6]), .A2(n247), .ZN(N159) );
  AND2_X1 U138 ( .A1(jump_address_dec[6]), .A2(n253), .ZN(N31) );
  AND2_X1 U139 ( .A1(immediate_dec[7]), .A2(n250), .ZN(N192) );
  AND2_X1 U140 ( .A1(immediate_ext_dec[7]), .A2(n247), .ZN(N160) );
  AND2_X1 U141 ( .A1(jump_address_dec[7]), .A2(n253), .ZN(N32) );
  AND2_X1 U142 ( .A1(immediate_dec[8]), .A2(n250), .ZN(N193) );
  AND2_X1 U143 ( .A1(immediate_ext_dec[8]), .A2(n247), .ZN(N161) );
  AND2_X1 U144 ( .A1(jump_address_dec[8]), .A2(n253), .ZN(N33) );
  AND2_X1 U145 ( .A1(immediate_dec[9]), .A2(n250), .ZN(N194) );
  AND2_X1 U146 ( .A1(immediate_ext_dec[9]), .A2(n247), .ZN(N162) );
  AND2_X1 U147 ( .A1(jump_address_dec[9]), .A2(n253), .ZN(N34) );
  AND2_X1 U148 ( .A1(immediate_dec[10]), .A2(n250), .ZN(N195) );
  AND2_X1 U149 ( .A1(immediate_ext_dec[10]), .A2(n247), .ZN(N163) );
  AND2_X1 U150 ( .A1(jump_address_dec[10]), .A2(n253), .ZN(N35) );
  AND2_X1 U151 ( .A1(rd_dec[0]), .A2(n251), .ZN(N206) );
  AND2_X1 U152 ( .A1(rd_dec[1]), .A2(n251), .ZN(N207) );
  AND2_X1 U153 ( .A1(rd_dec[2]), .A2(n251), .ZN(N208) );
  AND2_X1 U154 ( .A1(rd_dec[3]), .A2(n252), .ZN(N209) );
  AND2_X1 U155 ( .A1(immediate_dec[11]), .A2(n250), .ZN(N196) );
  AND2_X1 U156 ( .A1(immediate_dec[12]), .A2(n250), .ZN(N197) );
  AND2_X1 U157 ( .A1(immediate_dec[13]), .A2(n251), .ZN(N198) );
  AND2_X1 U158 ( .A1(immediate_dec[14]), .A2(n251), .ZN(N199) );
  AND2_X1 U159 ( .A1(immediate_ext_dec[11]), .A2(n247), .ZN(N164) );
  AND2_X1 U160 ( .A1(immediate_ext_dec[12]), .A2(n248), .ZN(N165) );
  AND2_X1 U161 ( .A1(immediate_ext_dec[13]), .A2(n248), .ZN(N166) );
  AND2_X1 U162 ( .A1(immediate_ext_dec[14]), .A2(n248), .ZN(N167) );
  AND2_X1 U163 ( .A1(read_data_1_dec[0]), .A2(n258), .ZN(N89) );
  AND2_X1 U164 ( .A1(read_data_1_dec[1]), .A2(n258), .ZN(N90) );
  AND2_X1 U165 ( .A1(read_data_1_dec[11]), .A2(n242), .ZN(N100) );
  AND2_X1 U166 ( .A1(read_data_1_dec[12]), .A2(n242), .ZN(N101) );
  AND2_X1 U167 ( .A1(read_data_1_dec[13]), .A2(n242), .ZN(N102) );
  AND2_X1 U168 ( .A1(read_data_1_dec[14]), .A2(n242), .ZN(N103) );
  AND2_X1 U169 ( .A1(read_data_1_dec[15]), .A2(n242), .ZN(N104) );
  AND2_X1 U170 ( .A1(read_data_1_dec[16]), .A2(n242), .ZN(N105) );
  AND2_X1 U171 ( .A1(read_data_1_dec[17]), .A2(n242), .ZN(N106) );
  AND2_X1 U172 ( .A1(read_data_1_dec[18]), .A2(n242), .ZN(N107) );
  AND2_X1 U173 ( .A1(read_data_1_dec[19]), .A2(n242), .ZN(N108) );
  AND2_X1 U174 ( .A1(read_data_1_dec[20]), .A2(n242), .ZN(N109) );
  AND2_X1 U175 ( .A1(read_data_1_dec[21]), .A2(n243), .ZN(N110) );
  AND2_X1 U176 ( .A1(read_data_1_dec[22]), .A2(n243), .ZN(N111) );
  AND2_X1 U177 ( .A1(read_data_1_dec[23]), .A2(n243), .ZN(N112) );
  AND2_X1 U178 ( .A1(read_data_1_dec[24]), .A2(n243), .ZN(N113) );
  AND2_X1 U179 ( .A1(read_data_1_dec[25]), .A2(n243), .ZN(N114) );
  AND2_X1 U180 ( .A1(read_data_1_dec[26]), .A2(n243), .ZN(N115) );
  AND2_X1 U181 ( .A1(read_data_1_dec[27]), .A2(n243), .ZN(N116) );
  AND2_X1 U182 ( .A1(read_data_1_dec[28]), .A2(n243), .ZN(N117) );
  AND2_X1 U183 ( .A1(read_data_1_dec[29]), .A2(n243), .ZN(N118) );
  AND2_X1 U184 ( .A1(read_data_1_dec[30]), .A2(n243), .ZN(N119) );
  AND2_X1 U185 ( .A1(read_data_1_dec[31]), .A2(n243), .ZN(N120) );
  AND2_X1 U186 ( .A1(pc_4_dec[0]), .A2(n255), .ZN(N57) );
  AND2_X1 U187 ( .A1(pc_4_dec[1]), .A2(n255), .ZN(N58) );
  AND2_X1 U188 ( .A1(pc_4_dec[2]), .A2(n256), .ZN(N59) );
  AND2_X1 U189 ( .A1(pc_4_dec[3]), .A2(n256), .ZN(N60) );
  AND2_X1 U190 ( .A1(pc_4_dec[4]), .A2(n256), .ZN(N61) );
  AND2_X1 U191 ( .A1(pc_4_dec[5]), .A2(n256), .ZN(N62) );
  AND2_X1 U192 ( .A1(pc_4_dec[6]), .A2(n256), .ZN(N63) );
  AND2_X1 U193 ( .A1(pc_4_dec[7]), .A2(n256), .ZN(N64) );
  AND2_X1 U194 ( .A1(pc_4_dec[8]), .A2(n256), .ZN(N65) );
  AND2_X1 U195 ( .A1(pc_4_dec[9]), .A2(n256), .ZN(N66) );
  AND2_X1 U196 ( .A1(pc_4_dec[10]), .A2(n256), .ZN(N67) );
  AND2_X1 U197 ( .A1(pc_4_dec[11]), .A2(n256), .ZN(N68) );
  AND2_X1 U198 ( .A1(pc_4_dec[12]), .A2(n256), .ZN(N69) );
  AND2_X1 U199 ( .A1(pc_4_dec[13]), .A2(n257), .ZN(N70) );
  AND2_X1 U200 ( .A1(pc_4_dec[14]), .A2(n257), .ZN(N71) );
  AND2_X1 U201 ( .A1(pc_4_dec[15]), .A2(n257), .ZN(N72) );
  AND2_X1 U202 ( .A1(pc_4_dec[16]), .A2(n257), .ZN(N73) );
  AND2_X1 U203 ( .A1(pc_4_dec[17]), .A2(n257), .ZN(N74) );
  AND2_X1 U204 ( .A1(pc_4_dec[18]), .A2(n257), .ZN(N75) );
  AND2_X1 U205 ( .A1(pc_4_dec[19]), .A2(n257), .ZN(N76) );
  AND2_X1 U206 ( .A1(pc_4_dec[20]), .A2(n257), .ZN(N77) );
  AND2_X1 U207 ( .A1(pc_4_dec[21]), .A2(n257), .ZN(N78) );
  AND2_X1 U208 ( .A1(pc_4_dec[22]), .A2(n257), .ZN(N79) );
  AND2_X1 U209 ( .A1(pc_4_dec[23]), .A2(n258), .ZN(N80) );
  AND2_X1 U210 ( .A1(pc_4_dec[24]), .A2(n258), .ZN(N81) );
  AND2_X1 U211 ( .A1(pc_4_dec[25]), .A2(n258), .ZN(N82) );
  AND2_X1 U212 ( .A1(pc_4_dec[26]), .A2(n258), .ZN(N83) );
  AND2_X1 U213 ( .A1(pc_4_dec[27]), .A2(n258), .ZN(N84) );
  AND2_X1 U214 ( .A1(pc_4_dec[28]), .A2(n258), .ZN(N85) );
  AND2_X1 U215 ( .A1(pc_4_dec[29]), .A2(n258), .ZN(N86) );
  AND2_X1 U216 ( .A1(pc_4_dec[30]), .A2(n258), .ZN(N87) );
  AND2_X1 U217 ( .A1(pc_4_dec[31]), .A2(n258), .ZN(N88) );
  AND2_X1 U218 ( .A1(jump_address_dec[11]), .A2(n253), .ZN(N36) );
  AND2_X1 U219 ( .A1(jump_address_dec[12]), .A2(n254), .ZN(N37) );
  AND2_X1 U220 ( .A1(jump_address_dec[13]), .A2(n254), .ZN(N38) );
  AND2_X1 U221 ( .A1(jump_address_dec[14]), .A2(n254), .ZN(N39) );
  AND2_X1 U222 ( .A1(cw_to_ex_dec[2]), .A2(n255), .ZN(N5) );
  AND2_X1 U223 ( .A1(cw_to_ex_dec[3]), .A2(n256), .ZN(N6) );
  AND2_X1 U224 ( .A1(cw_to_ex_dec[4]), .A2(n257), .ZN(N7) );
  AND2_X1 U225 ( .A1(cw_to_ex_dec[11]), .A2(n245), .ZN(N14) );
  AND2_X1 U226 ( .A1(cw_to_ex_dec[14]), .A2(n248), .ZN(N17) );
  AND2_X1 U227 ( .A1(cw_to_ex_dec[15]), .A2(n249), .ZN(N18) );
  AND2_X1 U228 ( .A1(cw_to_ex_dec[19]), .A2(n252), .ZN(N22) );
  AND2_X1 U229 ( .A1(read_data_1_dec[2]), .A2(n259), .ZN(N91) );
  AND2_X1 U230 ( .A1(read_data_1_dec[3]), .A2(n259), .ZN(N92) );
  AND2_X1 U231 ( .A1(read_data_1_dec[4]), .A2(n259), .ZN(N93) );
  AND2_X1 U232 ( .A1(read_data_1_dec[5]), .A2(n259), .ZN(N94) );
  AND2_X1 U233 ( .A1(read_data_1_dec[6]), .A2(n259), .ZN(N95) );
  AND2_X1 U234 ( .A1(read_data_1_dec[7]), .A2(n259), .ZN(N96) );
  AND2_X1 U235 ( .A1(read_data_1_dec[8]), .A2(n259), .ZN(N97) );
  AND2_X1 U236 ( .A1(read_data_1_dec[9]), .A2(n259), .ZN(N98) );
  AND2_X1 U237 ( .A1(read_data_1_dec[10]), .A2(n259), .ZN(N99) );
endmodule


module decode_unit ( address_write, data_write, pc_4_from_dec, instruction, 
        idex_rt, clk, rst, reg_write, idex_mem_read, cw, cw_to_ex, 
        jump_address, pc_4_to_ex, data_read_1, data_read_2, immediate_ext, 
        immediate, rt, rd, rs, opcode, func, pcwrite, ifid_write );
  input [4:0] address_write;
  input [31:0] data_write;
  input [31:0] pc_4_from_dec;
  input [31:0] instruction;
  input [4:0] idex_rt;
  input [3:0] idex_mem_read;
  input [22:0] cw;
  output [21:0] cw_to_ex;
  output [31:0] jump_address;
  output [31:0] pc_4_to_ex;
  output [31:0] data_read_1;
  output [31:0] data_read_2;
  output [31:0] immediate_ext;
  output [15:0] immediate;
  output [4:0] rt;
  output [4:0] rd;
  output [4:0] rs;
  output [5:0] opcode;
  output [10:0] func;
  input clk, rst, reg_write;
  output pcwrite, ifid_write;
  wire   \instruction[15] , \instruction[14] , \instruction[13] ,
         \instruction[12] , \instruction[11] , \instruction[20] ,
         \instruction[19] , \instruction[18] , \instruction[17] ,
         \instruction[16] , \instruction[25] , \instruction[24] ,
         \instruction[23] , \instruction[22] , \instruction[21] ,
         \instruction[31] , \instruction[30] , \instruction[29] ,
         \instruction[28] , \instruction[27] , \instruction[26] ,
         \instruction[10] , \instruction[9] , \instruction[8] ,
         \instruction[7] , \instruction[6] , \instruction[5] ,
         \instruction[4] , \instruction[3] , \instruction[2] ,
         \instruction[1] , \instruction[0] , \cw_i[21] , mux_op_i;
  assign pc_4_to_ex[31] = pc_4_from_dec[31];
  assign pc_4_to_ex[30] = pc_4_from_dec[30];
  assign pc_4_to_ex[29] = pc_4_from_dec[29];
  assign pc_4_to_ex[28] = pc_4_from_dec[28];
  assign pc_4_to_ex[27] = pc_4_from_dec[27];
  assign pc_4_to_ex[26] = pc_4_from_dec[26];
  assign pc_4_to_ex[25] = pc_4_from_dec[25];
  assign pc_4_to_ex[24] = pc_4_from_dec[24];
  assign pc_4_to_ex[23] = pc_4_from_dec[23];
  assign pc_4_to_ex[22] = pc_4_from_dec[22];
  assign pc_4_to_ex[21] = pc_4_from_dec[21];
  assign pc_4_to_ex[20] = pc_4_from_dec[20];
  assign pc_4_to_ex[19] = pc_4_from_dec[19];
  assign pc_4_to_ex[18] = pc_4_from_dec[18];
  assign pc_4_to_ex[17] = pc_4_from_dec[17];
  assign pc_4_to_ex[16] = pc_4_from_dec[16];
  assign pc_4_to_ex[15] = pc_4_from_dec[15];
  assign pc_4_to_ex[14] = pc_4_from_dec[14];
  assign pc_4_to_ex[13] = pc_4_from_dec[13];
  assign pc_4_to_ex[12] = pc_4_from_dec[12];
  assign pc_4_to_ex[11] = pc_4_from_dec[11];
  assign pc_4_to_ex[10] = pc_4_from_dec[10];
  assign pc_4_to_ex[9] = pc_4_from_dec[9];
  assign pc_4_to_ex[8] = pc_4_from_dec[8];
  assign pc_4_to_ex[7] = pc_4_from_dec[7];
  assign pc_4_to_ex[6] = pc_4_from_dec[6];
  assign pc_4_to_ex[5] = pc_4_from_dec[5];
  assign pc_4_to_ex[4] = pc_4_from_dec[4];
  assign pc_4_to_ex[3] = pc_4_from_dec[3];
  assign pc_4_to_ex[2] = pc_4_from_dec[2];
  assign pc_4_to_ex[1] = pc_4_from_dec[1];
  assign pc_4_to_ex[0] = pc_4_from_dec[0];
  assign immediate[15] = \instruction[15] ;
  assign rd[4] = \instruction[15] ;
  assign \instruction[15]  = instruction[15];
  assign immediate[14] = \instruction[14] ;
  assign rd[3] = \instruction[14] ;
  assign \instruction[14]  = instruction[14];
  assign immediate[13] = \instruction[13] ;
  assign rd[2] = \instruction[13] ;
  assign \instruction[13]  = instruction[13];
  assign immediate[12] = \instruction[12] ;
  assign rd[1] = \instruction[12] ;
  assign \instruction[12]  = instruction[12];
  assign immediate[11] = \instruction[11] ;
  assign rd[0] = \instruction[11] ;
  assign \instruction[11]  = instruction[11];
  assign rt[4] = \instruction[20] ;
  assign \instruction[20]  = instruction[20];
  assign rt[3] = \instruction[19] ;
  assign \instruction[19]  = instruction[19];
  assign rt[2] = \instruction[18] ;
  assign \instruction[18]  = instruction[18];
  assign rt[1] = \instruction[17] ;
  assign \instruction[17]  = instruction[17];
  assign rt[0] = \instruction[16] ;
  assign \instruction[16]  = instruction[16];
  assign rs[4] = \instruction[25] ;
  assign \instruction[25]  = instruction[25];
  assign rs[3] = \instruction[24] ;
  assign \instruction[24]  = instruction[24];
  assign rs[2] = \instruction[23] ;
  assign \instruction[23]  = instruction[23];
  assign rs[1] = \instruction[22] ;
  assign \instruction[22]  = instruction[22];
  assign rs[0] = \instruction[21] ;
  assign \instruction[21]  = instruction[21];
  assign opcode[5] = \instruction[31] ;
  assign \instruction[31]  = instruction[31];
  assign opcode[4] = \instruction[30] ;
  assign \instruction[30]  = instruction[30];
  assign opcode[3] = \instruction[29] ;
  assign \instruction[29]  = instruction[29];
  assign opcode[2] = \instruction[28] ;
  assign \instruction[28]  = instruction[28];
  assign opcode[1] = \instruction[27] ;
  assign \instruction[27]  = instruction[27];
  assign opcode[0] = \instruction[26] ;
  assign \instruction[26]  = instruction[26];
  assign immediate[10] = \instruction[10] ;
  assign func[10] = \instruction[10] ;
  assign \instruction[10]  = instruction[10];
  assign immediate[9] = \instruction[9] ;
  assign func[9] = \instruction[9] ;
  assign \instruction[9]  = instruction[9];
  assign immediate[8] = \instruction[8] ;
  assign func[8] = \instruction[8] ;
  assign \instruction[8]  = instruction[8];
  assign immediate[7] = \instruction[7] ;
  assign func[7] = \instruction[7] ;
  assign \instruction[7]  = instruction[7];
  assign immediate[6] = \instruction[6] ;
  assign func[6] = \instruction[6] ;
  assign \instruction[6]  = instruction[6];
  assign immediate[5] = \instruction[5] ;
  assign func[5] = \instruction[5] ;
  assign \instruction[5]  = instruction[5];
  assign immediate[4] = \instruction[4] ;
  assign func[4] = \instruction[4] ;
  assign \instruction[4]  = instruction[4];
  assign immediate[3] = \instruction[3] ;
  assign func[3] = \instruction[3] ;
  assign \instruction[3]  = instruction[3];
  assign immediate[2] = \instruction[2] ;
  assign func[2] = \instruction[2] ;
  assign \instruction[2]  = instruction[2];
  assign immediate[1] = \instruction[1] ;
  assign func[1] = \instruction[1] ;
  assign \instruction[1]  = instruction[1];
  assign immediate[0] = \instruction[0] ;
  assign func[0] = \instruction[0] ;
  assign \instruction[0]  = instruction[0];

  hdu hdu_0 ( .clk(clk), .rst(rst), .idex_mem_read(idex_mem_read), .idex_rt(
        idex_rt), .rs({\instruction[25] , \instruction[24] , \instruction[23] , 
        \instruction[22] , \instruction[21] }), .rt({\instruction[20] , 
        \instruction[19] , \instruction[18] , \instruction[17] , 
        \instruction[16] }), .pcwrite(pcwrite), .ifidwrite(ifid_write), 
        .mux_op(mux_op_i) );
  mux_stall mux_stall0 ( .cw_from_cu(cw), .mux_op(mux_op_i), .cw_from_mux({
        cw_to_ex[21], \cw_i[21] , cw_to_ex[20:0]}) );
  sign_extender sign_extender0 ( .immediate_jump({\instruction[25] , 
        \instruction[24] , \instruction[23] , \instruction[22] , 
        \instruction[21] , \instruction[20] , \instruction[19] , 
        \instruction[18] , \instruction[17] , \instruction[16] , 
        \instruction[15] , \instruction[14] , \instruction[13] , 
        \instruction[12] , \instruction[11] , \instruction[10] , 
        \instruction[9] , \instruction[8] , \instruction[7] , \instruction[6] , 
        \instruction[5] , \instruction[4] , \instruction[3] , \instruction[2] , 
        \instruction[1] , \instruction[0] }), .extended_jump(jump_address) );
  extender extender0 ( .immediate({\instruction[15] , \instruction[14] , 
        \instruction[13] , \instruction[12] , \instruction[11] , 
        \instruction[10] , \instruction[9] , \instruction[8] , 
        \instruction[7] , \instruction[6] , \instruction[5] , \instruction[4] , 
        \instruction[3] , \instruction[2] , \instruction[1] , \instruction[0] }), .unsigned_value(\cw_i[21] ), .extended(immediate_ext) );
  reg_file reg_file0 ( .read_address_1({\instruction[25] , \instruction[24] , 
        \instruction[23] , \instruction[22] , \instruction[21] }), 
        .read_address_2({\instruction[20] , \instruction[19] , 
        \instruction[18] , \instruction[17] , \instruction[16] }), 
        .write_address(address_write), .write_data(data_write), .reg_write(
        reg_write), .rst(rst), .data_reg_1(data_read_1), .data_reg_2(
        data_read_2) );
endmodule


module ifid_reg ( pc_4, instruction_fetch, flush, ifid_write, clk, rst, 
        instruction_decode, new_pc );
  input [31:0] pc_4;
  input [31:0] instruction_fetch;
  output [31:0] instruction_decode;
  output [31:0] new_pc;
  input flush, ifid_write, clk, rst;
  wire   n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n197,
         n202, n64, n65, n66, n67, n68, n196, n198, n199, n200, n201, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276;

  DFFR_X1 \instruction_decode_reg[31]  ( .D(n197), .CK(clk), .RN(n271), .Q(
        instruction_decode[31]), .QN(n132) );
  DFFS_X1 \instruction_decode_reg[30]  ( .D(n195), .CK(clk), .SN(n276), .Q(
        instruction_decode[30]), .QN(n131) );
  DFFR_X1 \instruction_decode_reg[29]  ( .D(n194), .CK(clk), .RN(n273), .Q(
        instruction_decode[29]), .QN(n130) );
  DFFS_X1 \instruction_decode_reg[28]  ( .D(n193), .CK(clk), .SN(n276), .Q(
        instruction_decode[28]), .QN(n129) );
  DFFR_X1 \instruction_decode_reg[27]  ( .D(n192), .CK(clk), .RN(n273), .Q(
        instruction_decode[27]), .QN(n128) );
  DFFS_X1 \instruction_decode_reg[26]  ( .D(n191), .CK(clk), .SN(n276), .Q(
        instruction_decode[26]), .QN(n127) );
  DFFR_X1 \instruction_decode_reg[25]  ( .D(n190), .CK(clk), .RN(n273), .Q(
        instruction_decode[25]), .QN(n126) );
  DFFR_X1 \instruction_decode_reg[24]  ( .D(n189), .CK(clk), .RN(n273), .Q(
        instruction_decode[24]), .QN(n125) );
  DFFR_X1 \instruction_decode_reg[23]  ( .D(n188), .CK(clk), .RN(n272), .Q(
        instruction_decode[23]), .QN(n124) );
  DFFR_X1 \instruction_decode_reg[22]  ( .D(n187), .CK(clk), .RN(n273), .Q(
        instruction_decode[22]), .QN(n123) );
  DFFR_X1 \instruction_decode_reg[21]  ( .D(n186), .CK(clk), .RN(n273), .Q(
        instruction_decode[21]), .QN(n122) );
  DFFR_X1 \instruction_decode_reg[20]  ( .D(n185), .CK(clk), .RN(n273), .Q(
        instruction_decode[20]), .QN(n121) );
  DFFR_X1 \instruction_decode_reg[19]  ( .D(n184), .CK(clk), .RN(n272), .Q(
        instruction_decode[19]), .QN(n120) );
  DFFR_X1 \instruction_decode_reg[18]  ( .D(n183), .CK(clk), .RN(n273), .Q(
        instruction_decode[18]), .QN(n119) );
  DFFR_X1 \instruction_decode_reg[17]  ( .D(n182), .CK(clk), .RN(n273), .Q(
        instruction_decode[17]), .QN(n118) );
  DFFR_X1 \instruction_decode_reg[16]  ( .D(n181), .CK(clk), .RN(n273), .Q(
        instruction_decode[16]), .QN(n117) );
  DFFR_X1 \instruction_decode_reg[15]  ( .D(n180), .CK(clk), .RN(n273), .Q(
        instruction_decode[15]), .QN(n116) );
  DFFR_X1 \instruction_decode_reg[14]  ( .D(n179), .CK(clk), .RN(n274), .Q(
        instruction_decode[14]), .QN(n115) );
  DFFR_X1 \instruction_decode_reg[13]  ( .D(n178), .CK(clk), .RN(n274), .Q(
        instruction_decode[13]), .QN(n114) );
  DFFR_X1 \instruction_decode_reg[12]  ( .D(n177), .CK(clk), .RN(n274), .Q(
        instruction_decode[12]), .QN(n113) );
  DFFR_X1 \instruction_decode_reg[11]  ( .D(n176), .CK(clk), .RN(n274), .Q(
        instruction_decode[11]), .QN(n112) );
  DFFR_X1 \instruction_decode_reg[10]  ( .D(n175), .CK(clk), .RN(n274), .Q(
        instruction_decode[10]), .QN(n111) );
  DFFR_X1 \instruction_decode_reg[9]  ( .D(n174), .CK(clk), .RN(n274), .Q(
        instruction_decode[9]), .QN(n110) );
  DFFR_X1 \instruction_decode_reg[8]  ( .D(n173), .CK(clk), .RN(n274), .Q(
        instruction_decode[8]), .QN(n109) );
  DFFR_X1 \instruction_decode_reg[7]  ( .D(n172), .CK(clk), .RN(n274), .Q(
        instruction_decode[7]), .QN(n108) );
  DFFR_X1 \instruction_decode_reg[6]  ( .D(n171), .CK(clk), .RN(n272), .Q(
        instruction_decode[6]), .QN(n107) );
  DFFR_X1 \instruction_decode_reg[5]  ( .D(n170), .CK(clk), .RN(n272), .Q(
        instruction_decode[5]), .QN(n106) );
  DFFR_X1 \instruction_decode_reg[4]  ( .D(n169), .CK(clk), .RN(n272), .Q(
        instruction_decode[4]), .QN(n105) );
  DFFR_X1 \instruction_decode_reg[3]  ( .D(n168), .CK(clk), .RN(n272), .Q(
        instruction_decode[3]), .QN(n104) );
  DFFR_X1 \instruction_decode_reg[2]  ( .D(n167), .CK(clk), .RN(n272), .Q(
        instruction_decode[2]), .QN(n103) );
  DFFR_X1 \instruction_decode_reg[1]  ( .D(n166), .CK(clk), .RN(n272), .Q(
        instruction_decode[1]), .QN(n102) );
  DFFR_X1 \instruction_decode_reg[0]  ( .D(n165), .CK(clk), .RN(n272), .Q(
        instruction_decode[0]), .QN(n101) );
  DFFR_X1 \new_pc_reg[31]  ( .D(n164), .CK(clk), .RN(n272), .Q(new_pc[31]), 
        .QN(n69) );
  DFFR_X1 \new_pc_reg[30]  ( .D(n163), .CK(clk), .RN(n272), .Q(new_pc[30]), 
        .QN(n70) );
  DFFR_X1 \new_pc_reg[29]  ( .D(n162), .CK(clk), .RN(n272), .Q(new_pc[29]), 
        .QN(n71) );
  DFFR_X1 \new_pc_reg[28]  ( .D(n161), .CK(clk), .RN(n274), .Q(new_pc[28]), 
        .QN(n72) );
  DFFR_X1 \new_pc_reg[27]  ( .D(n160), .CK(clk), .RN(n274), .Q(new_pc[27]), 
        .QN(n73) );
  DFFR_X1 \new_pc_reg[26]  ( .D(n159), .CK(clk), .RN(n275), .Q(new_pc[26]), 
        .QN(n74) );
  DFFR_X1 \new_pc_reg[25]  ( .D(n158), .CK(clk), .RN(n275), .Q(new_pc[25]), 
        .QN(n75) );
  DFFR_X1 \new_pc_reg[24]  ( .D(n157), .CK(clk), .RN(n274), .Q(new_pc[24]), 
        .QN(n76) );
  DFFR_X1 \new_pc_reg[23]  ( .D(n156), .CK(clk), .RN(n274), .Q(new_pc[23]), 
        .QN(n77) );
  DFFR_X1 \new_pc_reg[22]  ( .D(n155), .CK(clk), .RN(n275), .Q(new_pc[22]), 
        .QN(n78) );
  DFFR_X1 \new_pc_reg[21]  ( .D(n154), .CK(clk), .RN(n275), .Q(new_pc[21]), 
        .QN(n79) );
  DFFR_X1 \new_pc_reg[20]  ( .D(n153), .CK(clk), .RN(n275), .Q(new_pc[20]), 
        .QN(n80) );
  DFFR_X1 \new_pc_reg[19]  ( .D(n152), .CK(clk), .RN(n275), .Q(new_pc[19]), 
        .QN(n81) );
  DFFR_X1 \new_pc_reg[18]  ( .D(n151), .CK(clk), .RN(n275), .Q(new_pc[18]), 
        .QN(n82) );
  DFFR_X1 \new_pc_reg[17]  ( .D(n150), .CK(clk), .RN(n271), .Q(new_pc[17]), 
        .QN(n83) );
  DFFR_X1 \new_pc_reg[16]  ( .D(n149), .CK(clk), .RN(n271), .Q(new_pc[16]), 
        .QN(n84) );
  DFFR_X1 \new_pc_reg[15]  ( .D(n148), .CK(clk), .RN(n271), .Q(new_pc[15]), 
        .QN(n85) );
  DFFR_X1 \new_pc_reg[14]  ( .D(n147), .CK(clk), .RN(n271), .Q(new_pc[14]), 
        .QN(n86) );
  DFFR_X1 \new_pc_reg[13]  ( .D(n146), .CK(clk), .RN(n271), .Q(new_pc[13]), 
        .QN(n87) );
  DFFR_X1 \new_pc_reg[12]  ( .D(n145), .CK(clk), .RN(n271), .Q(new_pc[12]), 
        .QN(n88) );
  DFFR_X1 \new_pc_reg[11]  ( .D(n144), .CK(clk), .RN(n271), .Q(new_pc[11]), 
        .QN(n89) );
  DFFR_X1 \new_pc_reg[10]  ( .D(n143), .CK(clk), .RN(n271), .Q(new_pc[10]), 
        .QN(n90) );
  DFFR_X1 \new_pc_reg[9]  ( .D(n142), .CK(clk), .RN(n271), .Q(new_pc[9]), .QN(
        n91) );
  DFFR_X1 \new_pc_reg[8]  ( .D(n141), .CK(clk), .RN(n271), .Q(new_pc[8]), .QN(
        n92) );
  DFFR_X1 \new_pc_reg[7]  ( .D(n140), .CK(clk), .RN(n271), .Q(new_pc[7]), .QN(
        n93) );
  DFFR_X1 \new_pc_reg[6]  ( .D(n139), .CK(clk), .RN(n275), .Q(new_pc[6]), .QN(
        n94) );
  DFFR_X1 \new_pc_reg[5]  ( .D(n138), .CK(clk), .RN(n275), .Q(new_pc[5]), .QN(
        n95) );
  DFFR_X1 \new_pc_reg[4]  ( .D(n137), .CK(clk), .RN(n275), .Q(new_pc[4]), .QN(
        n96) );
  DFFR_X1 \new_pc_reg[3]  ( .D(n136), .CK(clk), .RN(n275), .Q(new_pc[3]), .QN(
        n97) );
  DFFR_X1 \new_pc_reg[2]  ( .D(n135), .CK(clk), .RN(n275), .Q(new_pc[2]), .QN(
        n98) );
  DFFR_X1 \new_pc_reg[1]  ( .D(n134), .CK(clk), .RN(n276), .Q(new_pc[1]), .QN(
        n99) );
  DFFR_X1 \new_pc_reg[0]  ( .D(n133), .CK(clk), .RN(n273), .Q(new_pc[0]), .QN(
        n100) );
  BUF_X1 U3 ( .A(n65), .Z(n261) );
  BUF_X1 U4 ( .A(n65), .Z(n262) );
  BUF_X1 U5 ( .A(n65), .Z(n263) );
  BUF_X1 U6 ( .A(n65), .Z(n264) );
  BUF_X1 U7 ( .A(n65), .Z(n260) );
  BUF_X1 U8 ( .A(n64), .Z(n269) );
  BUF_X1 U9 ( .A(n64), .Z(n268) );
  BUF_X1 U10 ( .A(n64), .Z(n265) );
  BUF_X1 U11 ( .A(n64), .Z(n266) );
  BUF_X1 U12 ( .A(n64), .Z(n267) );
  NAND2_X1 U13 ( .A1(n67), .A2(n265), .ZN(n65) );
  INV_X1 U14 ( .A(flush), .ZN(n202) );
  OAI22_X1 U15 ( .A1(n268), .A2(n80), .B1(n261), .B2(n239), .ZN(n153) );
  INV_X1 U16 ( .A(pc_4[20]), .ZN(n239) );
  OAI22_X1 U17 ( .A1(n268), .A2(n77), .B1(n261), .B2(n236), .ZN(n156) );
  INV_X1 U18 ( .A(pc_4[23]), .ZN(n236) );
  OAI22_X1 U19 ( .A1(n268), .A2(n76), .B1(n262), .B2(n235), .ZN(n157) );
  INV_X1 U20 ( .A(pc_4[24]), .ZN(n235) );
  OAI22_X1 U21 ( .A1(n268), .A2(n73), .B1(n262), .B2(n232), .ZN(n160) );
  INV_X1 U22 ( .A(pc_4[27]), .ZN(n232) );
  OAI22_X1 U23 ( .A1(n268), .A2(n72), .B1(n262), .B2(n231), .ZN(n161) );
  INV_X1 U24 ( .A(pc_4[28]), .ZN(n231) );
  OAI22_X1 U25 ( .A1(n268), .A2(n82), .B1(n261), .B2(n241), .ZN(n151) );
  INV_X1 U26 ( .A(pc_4[18]), .ZN(n241) );
  OAI22_X1 U27 ( .A1(n269), .A2(n81), .B1(n261), .B2(n240), .ZN(n152) );
  INV_X1 U28 ( .A(pc_4[19]), .ZN(n240) );
  OAI22_X1 U29 ( .A1(n268), .A2(n79), .B1(n261), .B2(n238), .ZN(n154) );
  INV_X1 U30 ( .A(pc_4[21]), .ZN(n238) );
  OAI22_X1 U31 ( .A1(n268), .A2(n78), .B1(n261), .B2(n237), .ZN(n155) );
  INV_X1 U32 ( .A(pc_4[22]), .ZN(n237) );
  OAI22_X1 U33 ( .A1(n268), .A2(n75), .B1(n262), .B2(n234), .ZN(n158) );
  INV_X1 U34 ( .A(pc_4[25]), .ZN(n234) );
  OAI22_X1 U35 ( .A1(n268), .A2(n74), .B1(n262), .B2(n233), .ZN(n159) );
  INV_X1 U36 ( .A(pc_4[26]), .ZN(n233) );
  OAI22_X1 U37 ( .A1(n268), .A2(n71), .B1(n262), .B2(n230), .ZN(n162) );
  INV_X1 U38 ( .A(pc_4[29]), .ZN(n230) );
  OAI22_X1 U39 ( .A1(n268), .A2(n70), .B1(n262), .B2(n229), .ZN(n163) );
  INV_X1 U40 ( .A(pc_4[30]), .ZN(n229) );
  OAI22_X1 U41 ( .A1(n268), .A2(n69), .B1(n262), .B2(n228), .ZN(n164) );
  INV_X1 U42 ( .A(pc_4[31]), .ZN(n228) );
  OAI22_X1 U43 ( .A1(n270), .A2(n100), .B1(n260), .B2(n259), .ZN(n133) );
  INV_X1 U44 ( .A(pc_4[0]), .ZN(n259) );
  OAI22_X1 U45 ( .A1(n270), .A2(n99), .B1(n260), .B2(n258), .ZN(n134) );
  INV_X1 U46 ( .A(pc_4[1]), .ZN(n258) );
  OAI22_X1 U47 ( .A1(n270), .A2(n98), .B1(n260), .B2(n257), .ZN(n135) );
  INV_X1 U48 ( .A(pc_4[2]), .ZN(n257) );
  OAI22_X1 U49 ( .A1(n270), .A2(n97), .B1(n260), .B2(n256), .ZN(n136) );
  INV_X1 U50 ( .A(pc_4[3]), .ZN(n256) );
  OAI22_X1 U51 ( .A1(n270), .A2(n96), .B1(n260), .B2(n255), .ZN(n137) );
  INV_X1 U52 ( .A(pc_4[4]), .ZN(n255) );
  OAI22_X1 U53 ( .A1(n270), .A2(n95), .B1(n260), .B2(n254), .ZN(n138) );
  INV_X1 U54 ( .A(pc_4[5]), .ZN(n254) );
  OAI22_X1 U55 ( .A1(n269), .A2(n88), .B1(n261), .B2(n247), .ZN(n145) );
  INV_X1 U56 ( .A(pc_4[12]), .ZN(n247) );
  OAI22_X1 U57 ( .A1(n269), .A2(n87), .B1(n261), .B2(n246), .ZN(n146) );
  INV_X1 U58 ( .A(pc_4[13]), .ZN(n246) );
  OAI22_X1 U59 ( .A1(n269), .A2(n86), .B1(n261), .B2(n245), .ZN(n147) );
  INV_X1 U60 ( .A(pc_4[14]), .ZN(n245) );
  OAI22_X1 U61 ( .A1(n269), .A2(n85), .B1(n261), .B2(n244), .ZN(n148) );
  INV_X1 U62 ( .A(pc_4[15]), .ZN(n244) );
  OAI22_X1 U63 ( .A1(n269), .A2(n84), .B1(n261), .B2(n243), .ZN(n149) );
  INV_X1 U64 ( .A(pc_4[16]), .ZN(n243) );
  OAI22_X1 U65 ( .A1(n101), .A2(n267), .B1(n262), .B2(n227), .ZN(n165) );
  INV_X1 U66 ( .A(instruction_fetch[0]), .ZN(n227) );
  OAI22_X1 U67 ( .A1(n102), .A2(n267), .B1(n262), .B2(n226), .ZN(n166) );
  INV_X1 U68 ( .A(instruction_fetch[1]), .ZN(n226) );
  OAI22_X1 U69 ( .A1(n103), .A2(n267), .B1(n262), .B2(n225), .ZN(n167) );
  INV_X1 U70 ( .A(instruction_fetch[2]), .ZN(n225) );
  OAI22_X1 U71 ( .A1(n104), .A2(n267), .B1(n262), .B2(n224), .ZN(n168) );
  INV_X1 U72 ( .A(instruction_fetch[3]), .ZN(n224) );
  OAI22_X1 U73 ( .A1(n105), .A2(n267), .B1(n263), .B2(n223), .ZN(n169) );
  INV_X1 U74 ( .A(instruction_fetch[4]), .ZN(n223) );
  OAI22_X1 U75 ( .A1(n106), .A2(n267), .B1(n263), .B2(n222), .ZN(n170) );
  INV_X1 U76 ( .A(instruction_fetch[5]), .ZN(n222) );
  OAI22_X1 U77 ( .A1(n107), .A2(n267), .B1(n263), .B2(n221), .ZN(n171) );
  INV_X1 U78 ( .A(instruction_fetch[6]), .ZN(n221) );
  OAI22_X1 U79 ( .A1(n108), .A2(n267), .B1(n263), .B2(n220), .ZN(n172) );
  INV_X1 U80 ( .A(instruction_fetch[7]), .ZN(n220) );
  OAI22_X1 U81 ( .A1(n109), .A2(n266), .B1(n263), .B2(n219), .ZN(n173) );
  INV_X1 U82 ( .A(instruction_fetch[8]), .ZN(n219) );
  OAI22_X1 U83 ( .A1(n110), .A2(n266), .B1(n263), .B2(n218), .ZN(n174) );
  INV_X1 U84 ( .A(instruction_fetch[9]), .ZN(n218) );
  OAI22_X1 U85 ( .A1(n111), .A2(n266), .B1(n263), .B2(n217), .ZN(n175) );
  INV_X1 U86 ( .A(instruction_fetch[10]), .ZN(n217) );
  OAI22_X1 U87 ( .A1(n112), .A2(n266), .B1(n263), .B2(n216), .ZN(n176) );
  INV_X1 U88 ( .A(instruction_fetch[11]), .ZN(n216) );
  OAI22_X1 U89 ( .A1(n113), .A2(n266), .B1(n263), .B2(n215), .ZN(n177) );
  INV_X1 U90 ( .A(instruction_fetch[12]), .ZN(n215) );
  OAI22_X1 U91 ( .A1(n114), .A2(n266), .B1(n263), .B2(n214), .ZN(n178) );
  INV_X1 U92 ( .A(instruction_fetch[13]), .ZN(n214) );
  OAI22_X1 U93 ( .A1(n115), .A2(n266), .B1(n263), .B2(n213), .ZN(n179) );
  INV_X1 U94 ( .A(instruction_fetch[14]), .ZN(n213) );
  OAI22_X1 U95 ( .A1(n116), .A2(n266), .B1(n263), .B2(n212), .ZN(n180) );
  INV_X1 U96 ( .A(instruction_fetch[15]), .ZN(n212) );
  OAI22_X1 U97 ( .A1(n117), .A2(n266), .B1(n264), .B2(n211), .ZN(n181) );
  INV_X1 U98 ( .A(instruction_fetch[16]), .ZN(n211) );
  OAI22_X1 U99 ( .A1(n118), .A2(n266), .B1(n264), .B2(n210), .ZN(n182) );
  INV_X1 U100 ( .A(instruction_fetch[17]), .ZN(n210) );
  OAI22_X1 U101 ( .A1(n119), .A2(n266), .B1(n264), .B2(n209), .ZN(n183) );
  INV_X1 U102 ( .A(instruction_fetch[18]), .ZN(n209) );
  OAI22_X1 U103 ( .A1(n120), .A2(n266), .B1(n264), .B2(n208), .ZN(n184) );
  INV_X1 U104 ( .A(instruction_fetch[19]), .ZN(n208) );
  OAI22_X1 U105 ( .A1(n121), .A2(n265), .B1(n264), .B2(n207), .ZN(n185) );
  INV_X1 U106 ( .A(instruction_fetch[20]), .ZN(n207) );
  OAI22_X1 U107 ( .A1(n122), .A2(n265), .B1(n264), .B2(n206), .ZN(n186) );
  INV_X1 U108 ( .A(instruction_fetch[21]), .ZN(n206) );
  OAI22_X1 U109 ( .A1(n123), .A2(n265), .B1(n264), .B2(n205), .ZN(n187) );
  INV_X1 U110 ( .A(instruction_fetch[22]), .ZN(n205) );
  OAI22_X1 U111 ( .A1(n124), .A2(n265), .B1(n264), .B2(n204), .ZN(n188) );
  INV_X1 U112 ( .A(instruction_fetch[23]), .ZN(n204) );
  OAI22_X1 U113 ( .A1(n125), .A2(n265), .B1(n264), .B2(n203), .ZN(n189) );
  INV_X1 U114 ( .A(instruction_fetch[24]), .ZN(n203) );
  OAI22_X1 U115 ( .A1(n126), .A2(n265), .B1(n264), .B2(n201), .ZN(n190) );
  INV_X1 U116 ( .A(instruction_fetch[25]), .ZN(n201) );
  OAI22_X1 U117 ( .A1(n128), .A2(n265), .B1(n264), .B2(n199), .ZN(n192) );
  INV_X1 U118 ( .A(instruction_fetch[27]), .ZN(n199) );
  OAI22_X1 U119 ( .A1(n130), .A2(n265), .B1(n264), .B2(n196), .ZN(n194) );
  INV_X1 U120 ( .A(instruction_fetch[29]), .ZN(n196) );
  OAI22_X1 U121 ( .A1(n269), .A2(n94), .B1(n260), .B2(n253), .ZN(n139) );
  INV_X1 U122 ( .A(pc_4[6]), .ZN(n253) );
  OAI22_X1 U123 ( .A1(n269), .A2(n93), .B1(n260), .B2(n252), .ZN(n140) );
  INV_X1 U124 ( .A(pc_4[7]), .ZN(n252) );
  OAI22_X1 U125 ( .A1(n269), .A2(n92), .B1(n260), .B2(n251), .ZN(n141) );
  INV_X1 U126 ( .A(pc_4[8]), .ZN(n251) );
  OAI22_X1 U127 ( .A1(n269), .A2(n91), .B1(n260), .B2(n250), .ZN(n142) );
  INV_X1 U128 ( .A(pc_4[9]), .ZN(n250) );
  OAI22_X1 U129 ( .A1(n269), .A2(n90), .B1(n260), .B2(n249), .ZN(n143) );
  INV_X1 U130 ( .A(pc_4[10]), .ZN(n249) );
  OAI22_X1 U131 ( .A1(n269), .A2(n89), .B1(n260), .B2(n248), .ZN(n144) );
  INV_X1 U132 ( .A(pc_4[11]), .ZN(n248) );
  OAI211_X1 U133 ( .C1(n127), .C2(n267), .A(n67), .B(n200), .ZN(n191) );
  NAND2_X1 U134 ( .A1(instruction_fetch[26]), .A2(n265), .ZN(n200) );
  OAI211_X1 U135 ( .C1(n129), .C2(n267), .A(n67), .B(n198), .ZN(n193) );
  NAND2_X1 U136 ( .A1(instruction_fetch[28]), .A2(n265), .ZN(n198) );
  OAI211_X1 U137 ( .C1(n131), .C2(n267), .A(n67), .B(n68), .ZN(n195) );
  NAND2_X1 U138 ( .A1(instruction_fetch[30]), .A2(n265), .ZN(n68) );
  INV_X1 U139 ( .A(rst), .ZN(n67) );
  OR2_X1 U140 ( .A1(ifid_write), .A2(rst), .ZN(n64) );
  OAI22_X1 U141 ( .A1(n132), .A2(n267), .B1(n65), .B2(n66), .ZN(n197) );
  INV_X1 U142 ( .A(instruction_fetch[31]), .ZN(n66) );
  OAI22_X1 U143 ( .A1(n269), .A2(n83), .B1(n261), .B2(n242), .ZN(n150) );
  INV_X1 U144 ( .A(pc_4[17]), .ZN(n242) );
  CLKBUF_X1 U145 ( .A(n64), .Z(n270) );
  CLKBUF_X1 U146 ( .A(n202), .Z(n271) );
  CLKBUF_X1 U147 ( .A(n202), .Z(n272) );
  CLKBUF_X1 U148 ( .A(n202), .Z(n273) );
  CLKBUF_X1 U149 ( .A(n202), .Z(n274) );
  CLKBUF_X1 U150 ( .A(n202), .Z(n275) );
  CLKBUF_X1 U151 ( .A(n202), .Z(n276) );
endmodule


module fetch ( jump_address, branch_target, from_iram, flush, clk, rst, pcsrc, 
        jump, pcwrite, to_iram, pc_4, instruction_fetch );
  input [31:0] jump_address;
  input [31:0] branch_target;
  input [31:0] from_iram;
  output [31:0] to_iram;
  output [31:0] pc_4;
  output [31:0] instruction_fetch;
  input flush, clk, rst, pcsrc, jump, pcwrite;

  wire   [31:0] data_mux_branch_i;
  wire   [31:0] data_mux_jump_i;
  wire   [31:0] data_pc_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign to_iram[31] = 1'b0;
  assign to_iram[30] = 1'b0;

  mux_branch mux_branch1 ( .from_increment_pc(pc_4), .branch_target(
        branch_target), .pcsrc(pcsrc), .to_mux_jump(data_mux_branch_i) );
  mux_jump mux_jump1 ( .jump_address(jump_address), .from_mux_branch(
        data_mux_branch_i), .jump(jump), .to_pc(data_mux_jump_i) );
  pc pc1 ( .from_mux_jump(data_mux_jump_i), .pcwrite(pcwrite), .clk(clk), 
        .rst(rst), .to_iram_block(data_pc_i) );
  increment_pc inc_pc1 ( .from_pc(data_pc_i), .to_mux_branch(pc_4) );
  iram_block iram_block1 ( .from_pc(data_pc_i), .flush(flush), .from_iram(
        from_iram), .to_iram({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        to_iram[29:0]}), .to_if_id_reg(instruction_fetch) );
endmodule


module DataPath ( clk, rst, fromIRAM, cw, Data_out_fromRAM, opcode, func, Addr, 
        read_op, write_op, nibble, write_byte, Address_toRAM, Data_in );
  input [31:0] fromIRAM;
  input [22:0] cw;
  input [31:0] Data_out_fromRAM;
  output [5:0] opcode;
  output [10:0] func;
  output [31:0] Addr;
  output [1:0] nibble;
  output [31:0] Address_toRAM;
  output [31:0] Data_in;
  input clk, rst;
  output read_op, write_op, write_byte;
  wire   flush_i, pcsrc_i, jump_i, pcwrite_i, ifid_write_i, reg_write_i,
         unaligned_i, regwriteMEM_i, branchTaken_i, takeBranch_out_i;
  wire   [31:0] jump_address_i;
  wire   [31:0] branch_target_i;
  wire   [31:0] pc_4_i;
  wire   [31:0] instruction_fetch_i;
  wire   [31:0] instruction_decode_i;
  wire   [31:0] new_pc_i;
  wire   [4:0] address_write_i;
  wire   [31:0] data_write_i;
  wire   [4:0] idex_rt_i;
  wire   [3:0] idex_mem_read_i;
  wire   [21:0] cw_to_idex_i;
  wire   [31:0] jaddr_i;
  wire   [31:0] pc4_to_idexreg_i;
  wire   [31:0] data_read_dec_1_i;
  wire   [31:0] data_read_dec_2_i;
  wire   [31:0] immediate_ext_dec_i;
  wire   [15:0] immediate_dec_i;
  wire   [4:0] rt_dec_i;
  wire   [4:0] rd_dec_i;
  wire   [4:0] rs_dec_i;
  wire   [21:0] cw_to_ex_i;
  wire   [31:0] jump_address_toex_i;
  wire   [31:0] pc_4_to_ex_i;
  wire   [31:0] data_read_ex_1_i;
  wire   [31:0] data_read_ex_2_i;
  wire   [31:0] immediate_ext_ex_i;
  wire   [15:0] immediate_ex_i;
  wire   [4:0] rt_ex_i;
  wire   [4:0] rd_ex_i;
  wire   [4:0] rs_ex_i;
  wire   [31:0] forw_dataMEM_i;
  wire   [4:0] RFaddr_MEM_i;
  wire   [10:0] cw_exmem_i;
  wire   [31:0] toPC1_i;
  wire   [31:0] toPC2_i;
  wire   [31:0] addrMem_exmem_i;
  wire   [31:0] writeData_exmem_i;
  wire   [4:0] addrRF_exmem_i;
  wire   [10:0] cw_tomem_i;
  wire   [31:0] PC1_tomem_i;
  wire   [31:0] PC2_tomem_i;
  wire   [31:0] mem_addr_out_i;
  wire   [31:0] mem_writedata_out_i;
  wire   [4:0] regfile_addr_out_tomem_i;
  wire   [2:0] cw_memwb_i;
  wire   [31:0] dataOut_mem_i;
  wire   [31:0] dataOut_exe_i;
  wire   [4:0] RFaddr_out_memwb_i;
  wire   [2:0] cw_towb_i;
  wire   [31:0] from_mem_data_out_i;
  wire   [31:0] from_alu_data_out_i;
  wire   [4:0] regfile_addr_out_towb_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign Addr[31] = 1'b0;
  assign Addr[30] = 1'b0;
  assign Address_toRAM[31] = 1'b0;
  assign Address_toRAM[30] = 1'b0;

  fetch u_fetch ( .jump_address(jump_address_i), .branch_target(
        branch_target_i), .from_iram(fromIRAM), .flush(flush_i), .clk(clk), 
        .rst(rst), .pcsrc(pcsrc_i), .jump(jump_i), .pcwrite(pcwrite_i), 
        .to_iram({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, Addr[29:0]}), .pc_4(pc_4_i), .instruction_fetch(instruction_fetch_i) );
  ifid_reg u_ifidreg ( .pc_4(pc_4_i), .instruction_fetch(instruction_fetch_i), 
        .flush(flush_i), .ifid_write(ifid_write_i), .clk(clk), .rst(rst), 
        .instruction_decode(instruction_decode_i), .new_pc(new_pc_i) );
  decode_unit u_decode_unit ( .address_write(address_write_i), .data_write(
        data_write_i), .pc_4_from_dec(new_pc_i), .instruction(
        instruction_decode_i), .idex_rt(idex_rt_i), .clk(clk), .rst(rst), 
        .reg_write(reg_write_i), .idex_mem_read(idex_mem_read_i), .cw(cw), 
        .cw_to_ex(cw_to_idex_i), .jump_address(jaddr_i), .pc_4_to_ex(
        pc4_to_idexreg_i), .data_read_1(data_read_dec_1_i), .data_read_2(
        data_read_dec_2_i), .immediate_ext(immediate_ext_dec_i), .immediate(
        immediate_dec_i), .rt(rt_dec_i), .rd(rd_dec_i), .rs(rs_dec_i), 
        .opcode(opcode), .func(func), .pcwrite(pcwrite_i), .ifid_write(
        ifid_write_i) );
  idex_reg u_idexreg ( .cw_to_ex_dec(cw_to_idex_i), .jump_address_dec(jaddr_i), 
        .pc_4_dec(pc4_to_idexreg_i), .read_data_1_dec(data_read_dec_1_i), 
        .read_data_2_dec(data_read_dec_2_i), .immediate_ext_dec(
        immediate_ext_dec_i), .immediate_dec(immediate_dec_i), .rt_dec(
        rt_dec_i), .rd_dec(rd_dec_i), .rs_dec(rs_dec_i), .clk(clk), .rst(rst), 
        .cw_to_ex(cw_to_ex_i), .jump_address(jump_address_toex_i), .pc_4(
        pc_4_to_ex_i), .read_data_1(data_read_ex_1_i), .read_data_2(
        data_read_ex_2_i), .immediate_ext(immediate_ext_ex_i), .immediate(
        immediate_ex_i), .rt(rt_ex_i), .rd(rd_ex_i), .rs(rs_ex_i) );
  execute u_execute ( .clk(clk), .rst(rst), .controls_in(cw_to_ex_i), 
        .ext25_0(jump_address_toex_i), .nextPC(pc_4_to_ex_i), .op_A(
        data_read_ex_1_i), .op_B(data_read_ex_2_i), .ext15_0(
        immediate_ext_ex_i), .inst15_0(immediate_ex_i), .rt_inst(rt_ex_i), 
        .rd_inst(rd_ex_i), .rs_inst(rs_ex_i), .unaligned(unaligned_i), 
        .forw_dataWB(data_write_i), .forw_dataMEM(forw_dataMEM_i), .RFaddr_WB(
        address_write_i), .RFaddr_MEM(RFaddr_MEM_i), .regwriteWB(reg_write_i), 
        .regwriteMEM(regwriteMEM_i), .controls_out(cw_exmem_i), .toPC1(toPC1_i), .toPC2(toPC2_i), .branchTaken(branchTaken_i), .addrMem(addrMem_exmem_i), 
        .writeData(writeData_exmem_i), .addrRF(addrRF_exmem_i), .IDEX_rt(
        idex_rt_i), .IDEX_memread(idex_mem_read_i) );
  EX_MEM_Reg u_exmemreg ( .clk(clk), .rst(rst), .controls_in(cw_exmem_i), 
        .toPC1_in(toPC1_i), .toPC2_in(toPC2_i), .takeBranch_in(branchTaken_i), 
        .mem_addr_in(addrMem_exmem_i), .mem_writedata_in(writeData_exmem_i), 
        .regfile_addr_in(addrRF_exmem_i), .controls_out(cw_tomem_i), 
        .toPC1_out(PC1_tomem_i), .toPC2_out(PC2_tomem_i), .takeBranch_out(
        takeBranch_out_i), .mem_addr_out(mem_addr_out_i), .mem_writedata_out(
        mem_writedata_out_i), .regfile_addr_out(regfile_addr_out_tomem_i) );
  memory u_memory ( .controls_in(cw_tomem_i), .PC1_in(PC1_tomem_i), .PC2_in(
        PC2_tomem_i), .takeBranch(takeBranch_out_i), .addrMem(mem_addr_out_i), 
        .writeData(mem_writedata_out_i), .RFaddr_in(regfile_addr_out_tomem_i), 
        .Data_out_fromRAM(Data_out_fromRAM), .controls_out(cw_memwb_i), 
        .dataOut_mem(dataOut_mem_i), .dataOut_exe(dataOut_exe_i), .RFaddr_out(
        RFaddr_out_memwb_i), .unaligned(unaligned_i), .PCsrc(pcsrc_i), .flush(
        flush_i), .jump(jump_i), .PC1_out(jump_address_i), .PC2_out(
        branch_target_i), .regwrite_MEM(regwriteMEM_i), .RFaddr_MEM(
        RFaddr_MEM_i), .forw_addr_MEM(forw_dataMEM_i), .read_op(read_op), 
        .write_op(write_op), .nibble(nibble), .write_byte(write_byte), 
        .Address_toRAM({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        Address_toRAM[29:0]}), .Data_in(Data_in) );
  MEM_WB_Reg u_memwbreg ( .clk(clk), .rst(rst), .controls_in(cw_memwb_i), 
        .from_mem_data_in(dataOut_mem_i), .from_alu_data_in(dataOut_exe_i), 
        .regfile_addr_in(RFaddr_out_memwb_i), .controls_out(cw_towb_i), 
        .from_mem_data_out(from_mem_data_out_i), .from_alu_data_out(
        from_alu_data_out_i), .regfile_addr_out(regfile_addr_out_towb_i) );
  writeback u_writeback ( .from_mem_data(from_mem_data_out_i), .from_alu_data(
        from_alu_data_out_i), .regfile_addr_in(regfile_addr_out_towb_i), 
        .regwrite_in(cw_towb_i[2]), .link(cw_towb_i[1]), .memtoreg(
        cw_towb_i[0]), .regwrite_out(reg_write_i), .regfile_data(data_write_i), 
        .regfile_addr_out(address_write_i) );
endmodule


module cu ( opcode, func, cw );
  input [5:0] opcode;
  input [10:0] func;
  output [22:0] cw;
  wire   n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  NAND3_X1 U115 ( .A1(cw[16]), .A2(n40), .A3(func[3]), .ZN(n36) );
  NAND3_X1 U116 ( .A1(opcode[1]), .A2(n45), .A3(n46), .ZN(n35) );
  NAND3_X1 U117 ( .A1(n81), .A2(n82), .A3(n83), .ZN(cw[1]) );
  XOR2_X1 U118 ( .A(func[1]), .B(n118), .Z(n117) );
  NAND3_X1 U119 ( .A1(opcode[4]), .A2(n45), .A3(n38), .ZN(n48) );
  NAND3_X1 U120 ( .A1(n30), .A2(n45), .A3(opcode[1]), .ZN(n32) );
  NAND3_X1 U121 ( .A1(opcode[0]), .A2(n45), .A3(opcode[1]), .ZN(n79) );
  NAND3_X1 U122 ( .A1(func[5]), .A2(n43), .A3(func[1]), .ZN(n42) );
  NAND3_X1 U123 ( .A1(opcode[0]), .A2(n39), .A3(n46), .ZN(n107) );
  NAND3_X1 U124 ( .A1(func[3]), .A2(n118), .A3(n59), .ZN(n56) );
  INV_X1 U3 ( .A(n76), .ZN(n52) );
  INV_X1 U4 ( .A(n101), .ZN(n77) );
  INV_X1 U5 ( .A(cw[16]), .ZN(n120) );
  INV_X1 U6 ( .A(n109), .ZN(n80) );
  INV_X1 U7 ( .A(cw[18]), .ZN(n33) );
  INV_X1 U8 ( .A(n98), .ZN(n87) );
  INV_X1 U9 ( .A(n110), .ZN(n29) );
  INV_X1 U10 ( .A(n90), .ZN(n53) );
  INV_X1 U11 ( .A(cw[12]), .ZN(n100) );
  NOR2_X1 U12 ( .A1(n31), .A2(n101), .ZN(cw[16]) );
  NOR3_X1 U13 ( .A1(n60), .A2(n120), .A3(n42), .ZN(n73) );
  AOI211_X1 U14 ( .C1(cw[16]), .C2(n124), .A(n47), .B(n66), .ZN(n82) );
  NAND4_X1 U15 ( .A1(n30), .A2(n91), .A3(n45), .A4(n123), .ZN(n101) );
  OAI22_X1 U16 ( .A1(n79), .A2(n108), .B1(n80), .B2(n94), .ZN(n92) );
  INV_X1 U17 ( .A(n46), .ZN(n108) );
  OAI22_X1 U18 ( .A1(n79), .A2(n80), .B1(n93), .B2(n31), .ZN(cw[18]) );
  NOR2_X1 U19 ( .A1(n111), .A2(n123), .ZN(n46) );
  NOR2_X1 U20 ( .A1(n78), .A2(n62), .ZN(n110) );
  NAND2_X1 U21 ( .A1(n38), .A2(n123), .ZN(n76) );
  INV_X1 U22 ( .A(n85), .ZN(n38) );
  NOR2_X1 U23 ( .A1(n123), .A2(n31), .ZN(n109) );
  INV_X1 U24 ( .A(n119), .ZN(n39) );
  NAND2_X1 U25 ( .A1(cw[16]), .A2(n60), .ZN(n98) );
  NOR2_X1 U26 ( .A1(n111), .A2(n93), .ZN(cw[12]) );
  NAND2_X1 U27 ( .A1(n101), .A2(n93), .ZN(n68) );
  NAND2_X1 U28 ( .A1(n73), .A2(n41), .ZN(n50) );
  NAND2_X1 U29 ( .A1(n52), .A2(n30), .ZN(n90) );
  INV_X1 U30 ( .A(n56), .ZN(n124) );
  OR3_X1 U31 ( .A1(cw[10]), .A2(cw[8]), .A3(n110), .ZN(cw[7]) );
  NAND4_X1 U32 ( .A1(n104), .A2(n105), .A3(n106), .A4(n107), .ZN(cw[21]) );
  INV_X1 U33 ( .A(n92), .ZN(n104) );
  NAND2_X1 U34 ( .A1(n52), .A2(n69), .ZN(n106) );
  AOI211_X1 U35 ( .C1(n39), .C2(n38), .A(n102), .B(n103), .ZN(n74) );
  INV_X1 U36 ( .A(n48), .ZN(n102) );
  OR2_X1 U37 ( .A1(cw[7]), .A2(cw[21]), .ZN(n103) );
  INV_X1 U38 ( .A(n47), .ZN(n34) );
  NAND4_X1 U39 ( .A1(n82), .A2(n105), .A3(n112), .A4(n113), .ZN(cw[0]) );
  NOR4_X1 U40 ( .A1(n110), .A2(n71), .A3(n114), .A4(n115), .ZN(n113) );
  AOI21_X1 U41 ( .B1(n71), .B2(n91), .A(n92), .ZN(n81) );
  OAI21_X1 U42 ( .B1(n31), .B2(n32), .A(n33), .ZN(cw[6]) );
  NOR2_X1 U43 ( .A1(n29), .A2(n30), .ZN(cw[9]) );
  NOR2_X1 U44 ( .A1(n101), .A2(n111), .ZN(cw[13]) );
  NOR3_X1 U45 ( .A1(n94), .A2(n30), .A3(n76), .ZN(cw[17]) );
  AOI21_X1 U46 ( .B1(n79), .B2(n32), .A(n80), .ZN(cw[20]) );
  NAND4_X1 U47 ( .A1(n74), .A2(n75), .A3(n76), .A4(n33), .ZN(cw[22]) );
  NAND2_X1 U48 ( .A1(n77), .A2(n78), .ZN(n75) );
  NOR4_X1 U49 ( .A1(n89), .A2(n41), .A3(n118), .A4(func[1]), .ZN(n95) );
  OAI221_X1 U50 ( .B1(n125), .B2(n120), .C1(n79), .C2(n76), .A(n49), .ZN(n66)
         );
  AOI21_X1 U51 ( .B1(n124), .B2(func[2]), .A(n126), .ZN(n125) );
  NOR4_X1 U52 ( .A1(func[4]), .A2(func[3]), .A3(n118), .A4(n42), .ZN(n126) );
  NOR4_X1 U53 ( .A1(func[9]), .A2(func[8]), .A3(func[7]), .A4(func[6]), .ZN(
        n97) );
  INV_X1 U54 ( .A(opcode[0]), .ZN(n30) );
  AOI211_X1 U55 ( .C1(n52), .C2(n45), .A(n65), .B(n66), .ZN(n64) );
  INV_X1 U56 ( .A(n67), .ZN(n65) );
  AOI22_X1 U57 ( .A1(n68), .A2(opcode[5]), .B1(n69), .B2(n38), .ZN(n67) );
  NOR3_X1 U58 ( .A1(n78), .A2(opcode[3]), .A3(n101), .ZN(cw[8]) );
  NOR3_X1 U59 ( .A1(n78), .A2(opcode[3]), .A3(n93), .ZN(cw[10]) );
  NOR2_X1 U60 ( .A1(n48), .A2(opcode[0]), .ZN(n71) );
  AOI22_X1 U61 ( .A1(n121), .A2(n46), .B1(n122), .B2(n109), .ZN(n105) );
  INV_X1 U62 ( .A(n32), .ZN(n121) );
  OAI22_X1 U63 ( .A1(n94), .A2(n30), .B1(n119), .B2(opcode[0]), .ZN(n122) );
  NOR3_X1 U64 ( .A1(n76), .A2(opcode[1]), .A3(n30), .ZN(n114) );
  INV_X1 U65 ( .A(func[4]), .ZN(n41) );
  NOR2_X1 U66 ( .A1(n61), .A2(func[1]), .ZN(n59) );
  OAI22_X1 U67 ( .A1(n41), .A2(n42), .B1(n43), .B2(n44), .ZN(n40) );
  NAND4_X1 U68 ( .A1(n38), .A2(opcode[4]), .A3(n39), .A4(n30), .ZN(n49) );
  AOI22_X1 U69 ( .A1(n73), .A2(n118), .B1(opcode[5]), .B2(n68), .ZN(n112) );
  NOR2_X1 U70 ( .A1(n30), .A2(opcode[2]), .ZN(n69) );
  INV_X1 U71 ( .A(opcode[5]), .ZN(n78) );
  NAND2_X1 U72 ( .A1(opcode[1]), .A2(opcode[2]), .ZN(n94) );
  INV_X1 U73 ( .A(func[0]), .ZN(n118) );
  AOI21_X1 U74 ( .B1(n44), .B2(n116), .A(n98), .ZN(n115) );
  NAND4_X1 U75 ( .A1(n117), .A2(func[2]), .A3(n41), .A4(n89), .ZN(n116) );
  NAND2_X1 U76 ( .A1(n59), .A2(func[0]), .ZN(n44) );
  NAND2_X1 U77 ( .A1(opcode[3]), .A2(opcode[5]), .ZN(n111) );
  INV_X1 U78 ( .A(func[2]), .ZN(n43) );
  AOI21_X1 U79 ( .B1(n44), .B2(n72), .A(func[2]), .ZN(n70) );
  OR2_X1 U80 ( .A1(n61), .A2(func[3]), .ZN(n72) );
  OAI211_X1 U81 ( .C1(n44), .C2(n55), .A(n56), .B(n57), .ZN(n54) );
  NAND2_X1 U82 ( .A1(func[3]), .A2(n43), .ZN(n55) );
  OAI211_X1 U83 ( .C1(n58), .C2(n59), .A(n60), .B(func[2]), .ZN(n57) );
  NOR2_X1 U84 ( .A1(func[0]), .A2(n61), .ZN(n58) );
  INV_X1 U85 ( .A(opcode[2]), .ZN(n45) );
  AOI221_X1 U86 ( .B1(n73), .B2(func[0]), .C1(n53), .C2(opcode[1]), .A(n84), 
        .ZN(n83) );
  OAI21_X1 U87 ( .B1(n79), .B2(n85), .A(n86), .ZN(n84) );
  NAND4_X1 U88 ( .A1(n87), .A2(func[1]), .A3(n88), .A4(n41), .ZN(n86) );
  OAI22_X1 U89 ( .A1(func[5]), .A2(n43), .B1(func[0]), .B2(n89), .ZN(n88) );
  NAND4_X1 U90 ( .A1(n38), .A2(opcode[4]), .A3(opcode[0]), .A4(n39), .ZN(n37)
         );
  INV_X1 U91 ( .A(opcode[4]), .ZN(n123) );
  OR2_X1 U92 ( .A1(n79), .A2(opcode[4]), .ZN(n93) );
  OR2_X1 U93 ( .A1(opcode[3]), .A2(opcode[5]), .ZN(n31) );
  NAND2_X1 U94 ( .A1(opcode[3]), .A2(n78), .ZN(n85) );
  NAND2_X1 U95 ( .A1(opcode[2]), .A2(n91), .ZN(n119) );
  NAND2_X1 U96 ( .A1(func[5]), .A2(n41), .ZN(n61) );
  INV_X1 U97 ( .A(func[3]), .ZN(n60) );
  INV_X1 U98 ( .A(opcode[1]), .ZN(n91) );
  NOR2_X1 U99 ( .A1(n62), .A2(opcode[5]), .ZN(cw[5]) );
  INV_X1 U100 ( .A(func[5]), .ZN(n89) );
  NAND2_X1 U101 ( .A1(n107), .A2(n127), .ZN(n47) );
  NAND4_X1 U102 ( .A1(func[3]), .A2(func[2]), .A3(cw[16]), .A4(n95), .ZN(n127)
         );
  OR3_X1 U103 ( .A1(opcode[3]), .A2(opcode[4]), .A3(n119), .ZN(n62) );
  NAND4_X1 U104 ( .A1(n50), .A2(n62), .A3(n63), .A4(n64), .ZN(cw[2]) );
  AOI22_X1 U105 ( .A1(n70), .A2(cw[16]), .B1(n71), .B2(opcode[1]), .ZN(n63) );
  NAND4_X1 U106 ( .A1(n48), .A2(n49), .A3(n50), .A4(n51), .ZN(cw[3]) );
  AOI222_X1 U107 ( .A1(n52), .A2(n39), .B1(n53), .B2(opcode[2]), .C1(cw[16]), 
        .C2(n54), .ZN(n51) );
  NAND4_X1 U108 ( .A1(n34), .A2(n35), .A3(n36), .A4(n37), .ZN(cw[4]) );
  NOR2_X1 U109 ( .A1(opcode[0]), .A2(n29), .ZN(cw[11]) );
  NAND4_X1 U110 ( .A1(n74), .A2(n99), .A3(n90), .A4(n100), .ZN(cw[14]) );
  NAND2_X1 U111 ( .A1(opcode[3]), .A2(n77), .ZN(n99) );
  AND4_X1 U112 ( .A1(n87), .A2(n95), .A3(n96), .A4(n97), .ZN(cw[15]) );
  NOR2_X1 U113 ( .A1(func[2]), .A2(func[10]), .ZN(n96) );
  AND2_X1 U114 ( .A1(opcode[0]), .A2(cw[5]), .ZN(cw[19]) );
endmodule


module DLX ( clk, rst, iram_data, Data_out_fromRAM, addr_to_iram, read_op, 
        write_op, nibble, write_byte, Address_toRAM, Data_in );
  input [31:0] iram_data;
  input [31:0] Data_out_fromRAM;
  output [31:0] addr_to_iram;
  output [1:0] nibble;
  output [31:0] Address_toRAM;
  output [31:0] Data_in;
  input clk, rst;
  output read_op, write_op, write_byte;

  wire   [5:0] opcode_i;
  wire   [10:0] func_i;
  wire   [22:0] cw_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign addr_to_iram[31] = 1'b0;
  assign addr_to_iram[30] = 1'b0;
  assign Address_toRAM[31] = 1'b0;
  assign Address_toRAM[30] = 1'b0;

  cu u_cu ( .opcode(opcode_i), .func(func_i), .cw(cw_i) );
  DataPath u_DataPath ( .clk(clk), .rst(rst), .fromIRAM(iram_data), .cw(cw_i), 
        .Data_out_fromRAM(Data_out_fromRAM), .opcode(opcode_i), .func(func_i), 
        .Addr({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        addr_to_iram[29:0]}), .read_op(read_op), .write_op(write_op), .nibble(
        nibble), .write_byte(write_byte), .Address_toRAM({
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, Address_toRAM[29:0]}), .Data_in(Data_in) );
endmodule

